magic
tech sky130A
magscale 1 2
timestamp 1709561889
<< error_p >>
rect -147 281 -89 287
rect -29 281 29 287
rect 89 281 147 287
rect -147 247 -135 281
rect -29 247 -17 281
rect 89 247 101 281
rect -147 241 -89 247
rect -29 241 29 247
rect 89 241 147 247
rect -147 -247 -89 -241
rect -29 -247 29 -241
rect 89 -247 147 -241
rect -147 -281 -135 -247
rect -29 -281 -17 -247
rect 89 -281 101 -247
rect -147 -287 -89 -281
rect -29 -287 29 -281
rect 89 -287 147 -281
<< nwell >>
rect -344 -419 344 419
<< pmos >>
rect -148 -200 -88 200
rect -30 -200 30 200
rect 88 -200 148 200
<< pdiff >>
rect -206 188 -148 200
rect -206 -188 -194 188
rect -160 -188 -148 188
rect -206 -200 -148 -188
rect -88 188 -30 200
rect -88 -188 -76 188
rect -42 -188 -30 188
rect -88 -200 -30 -188
rect 30 188 88 200
rect 30 -188 42 188
rect 76 -188 88 188
rect 30 -200 88 -188
rect 148 188 206 200
rect 148 -188 160 188
rect 194 -188 206 188
rect 148 -200 206 -188
<< pdiffc >>
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
<< nsubdiff >>
rect -308 349 -212 383
rect 212 349 308 383
rect -308 287 -274 349
rect 274 287 308 349
rect -308 -349 -274 -287
rect 274 -349 308 -287
rect -308 -383 -212 -349
rect 212 -383 308 -349
<< nsubdiffcont >>
rect -212 349 212 383
rect -308 -287 -274 287
rect 274 -287 308 287
rect -212 -383 212 -349
<< poly >>
rect -151 281 -85 297
rect -151 247 -135 281
rect -101 247 -85 281
rect -151 231 -85 247
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect 85 281 151 297
rect 85 247 101 281
rect 135 247 151 281
rect 85 231 151 247
rect -148 200 -88 231
rect -30 200 30 231
rect 88 200 148 231
rect -148 -231 -88 -200
rect -30 -231 30 -200
rect 88 -231 148 -200
rect -151 -247 -85 -231
rect -151 -281 -135 -247
rect -101 -281 -85 -247
rect -151 -297 -85 -281
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
rect 85 -247 151 -231
rect 85 -281 101 -247
rect 135 -281 151 -247
rect 85 -297 151 -281
<< polycont >>
rect -135 247 -101 281
rect -17 247 17 281
rect 101 247 135 281
rect -135 -281 -101 -247
rect -17 -281 17 -247
rect 101 -281 135 -247
<< locali >>
rect -308 349 -212 383
rect 212 349 308 383
rect -308 287 -274 349
rect 274 287 308 349
rect -151 247 -135 281
rect -101 247 -85 281
rect -33 247 -17 281
rect 17 247 33 281
rect 85 247 101 281
rect 135 247 151 281
rect -194 188 -160 204
rect -194 -204 -160 -188
rect -76 188 -42 204
rect -76 -204 -42 -188
rect 42 188 76 204
rect 42 -204 76 -188
rect 160 188 194 204
rect 160 -204 194 -188
rect -151 -281 -135 -247
rect -101 -281 -85 -247
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect 85 -281 101 -247
rect 135 -281 151 -247
rect -308 -349 -274 -287
rect 274 -349 308 -287
rect -308 -383 -212 -349
rect 212 -383 308 -349
<< viali >>
rect -135 247 -101 281
rect -17 247 17 281
rect 101 247 135 281
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect -135 -281 -101 -247
rect -17 -281 17 -247
rect 101 -281 135 -247
<< metal1 >>
rect -147 281 -89 287
rect -147 247 -135 281
rect -101 247 -89 281
rect -147 241 -89 247
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect 89 281 147 287
rect 89 247 101 281
rect 135 247 147 281
rect 89 241 147 247
rect -200 188 -154 200
rect -200 -188 -194 188
rect -160 -188 -154 188
rect -200 -200 -154 -188
rect -82 188 -36 200
rect -82 -188 -76 188
rect -42 -188 -36 188
rect -82 -200 -36 -188
rect 36 188 82 200
rect 36 -188 42 188
rect 76 -188 82 188
rect 36 -200 82 -188
rect 154 188 200 200
rect 154 -188 160 188
rect 194 -188 200 188
rect 154 -200 200 -188
rect -147 -247 -89 -241
rect -147 -281 -135 -247
rect -101 -281 -89 -247
rect -147 -287 -89 -281
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
rect 89 -247 147 -241
rect 89 -281 101 -247
rect 135 -281 147 -247
rect 89 -287 147 -281
<< properties >>
string FIXED_BBOX -291 -366 291 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 0.3 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
