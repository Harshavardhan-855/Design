magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< pwell >>
rect -1057 -310 1057 310
<< nmos >>
rect -861 -100 -741 100
rect -683 -100 -563 100
rect -505 -100 -385 100
rect -327 -100 -207 100
rect -149 -100 -29 100
rect 29 -100 149 100
rect 207 -100 327 100
rect 385 -100 505 100
rect 563 -100 683 100
rect 741 -100 861 100
<< ndiff >>
rect -919 88 -861 100
rect -919 -88 -907 88
rect -873 -88 -861 88
rect -919 -100 -861 -88
rect -741 88 -683 100
rect -741 -88 -729 88
rect -695 -88 -683 88
rect -741 -100 -683 -88
rect -563 88 -505 100
rect -563 -88 -551 88
rect -517 -88 -505 88
rect -563 -100 -505 -88
rect -385 88 -327 100
rect -385 -88 -373 88
rect -339 -88 -327 88
rect -385 -100 -327 -88
rect -207 88 -149 100
rect -207 -88 -195 88
rect -161 -88 -149 88
rect -207 -100 -149 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 149 88 207 100
rect 149 -88 161 88
rect 195 -88 207 88
rect 149 -100 207 -88
rect 327 88 385 100
rect 327 -88 339 88
rect 373 -88 385 88
rect 327 -100 385 -88
rect 505 88 563 100
rect 505 -88 517 88
rect 551 -88 563 88
rect 505 -100 563 -88
rect 683 88 741 100
rect 683 -88 695 88
rect 729 -88 741 88
rect 683 -100 741 -88
rect 861 88 919 100
rect 861 -88 873 88
rect 907 -88 919 88
rect 861 -100 919 -88
<< ndiffc >>
rect -907 -88 -873 88
rect -729 -88 -695 88
rect -551 -88 -517 88
rect -373 -88 -339 88
rect -195 -88 -161 88
rect -17 -88 17 88
rect 161 -88 195 88
rect 339 -88 373 88
rect 517 -88 551 88
rect 695 -88 729 88
rect 873 -88 907 88
<< psubdiff >>
rect -1021 240 -925 274
rect 925 240 1021 274
rect -1021 178 -987 240
rect 987 178 1021 240
rect -1021 -240 -987 -178
rect 987 -240 1021 -178
rect -1021 -274 -925 -240
rect 925 -274 1021 -240
<< psubdiffcont >>
rect -925 240 925 274
rect -1021 -178 -987 178
rect 987 -178 1021 178
rect -925 -274 925 -240
<< poly >>
rect -861 172 -741 188
rect -861 138 -845 172
rect -757 138 -741 172
rect -861 100 -741 138
rect -683 172 -563 188
rect -683 138 -667 172
rect -579 138 -563 172
rect -683 100 -563 138
rect -505 172 -385 188
rect -505 138 -489 172
rect -401 138 -385 172
rect -505 100 -385 138
rect -327 172 -207 188
rect -327 138 -311 172
rect -223 138 -207 172
rect -327 100 -207 138
rect -149 172 -29 188
rect -149 138 -133 172
rect -45 138 -29 172
rect -149 100 -29 138
rect 29 172 149 188
rect 29 138 45 172
rect 133 138 149 172
rect 29 100 149 138
rect 207 172 327 188
rect 207 138 223 172
rect 311 138 327 172
rect 207 100 327 138
rect 385 172 505 188
rect 385 138 401 172
rect 489 138 505 172
rect 385 100 505 138
rect 563 172 683 188
rect 563 138 579 172
rect 667 138 683 172
rect 563 100 683 138
rect 741 172 861 188
rect 741 138 757 172
rect 845 138 861 172
rect 741 100 861 138
rect -861 -138 -741 -100
rect -861 -172 -845 -138
rect -757 -172 -741 -138
rect -861 -188 -741 -172
rect -683 -138 -563 -100
rect -683 -172 -667 -138
rect -579 -172 -563 -138
rect -683 -188 -563 -172
rect -505 -138 -385 -100
rect -505 -172 -489 -138
rect -401 -172 -385 -138
rect -505 -188 -385 -172
rect -327 -138 -207 -100
rect -327 -172 -311 -138
rect -223 -172 -207 -138
rect -327 -188 -207 -172
rect -149 -138 -29 -100
rect -149 -172 -133 -138
rect -45 -172 -29 -138
rect -149 -188 -29 -172
rect 29 -138 149 -100
rect 29 -172 45 -138
rect 133 -172 149 -138
rect 29 -188 149 -172
rect 207 -138 327 -100
rect 207 -172 223 -138
rect 311 -172 327 -138
rect 207 -188 327 -172
rect 385 -138 505 -100
rect 385 -172 401 -138
rect 489 -172 505 -138
rect 385 -188 505 -172
rect 563 -138 683 -100
rect 563 -172 579 -138
rect 667 -172 683 -138
rect 563 -188 683 -172
rect 741 -138 861 -100
rect 741 -172 757 -138
rect 845 -172 861 -138
rect 741 -188 861 -172
<< polycont >>
rect -845 138 -757 172
rect -667 138 -579 172
rect -489 138 -401 172
rect -311 138 -223 172
rect -133 138 -45 172
rect 45 138 133 172
rect 223 138 311 172
rect 401 138 489 172
rect 579 138 667 172
rect 757 138 845 172
rect -845 -172 -757 -138
rect -667 -172 -579 -138
rect -489 -172 -401 -138
rect -311 -172 -223 -138
rect -133 -172 -45 -138
rect 45 -172 133 -138
rect 223 -172 311 -138
rect 401 -172 489 -138
rect 579 -172 667 -138
rect 757 -172 845 -138
<< locali >>
rect -1021 240 -925 274
rect 925 240 1021 274
rect -1021 178 -987 240
rect 987 178 1021 240
rect -861 138 -845 172
rect -757 138 -741 172
rect -683 138 -667 172
rect -579 138 -563 172
rect -505 138 -489 172
rect -401 138 -385 172
rect -327 138 -311 172
rect -223 138 -207 172
rect -149 138 -133 172
rect -45 138 -29 172
rect 29 138 45 172
rect 133 138 149 172
rect 207 138 223 172
rect 311 138 327 172
rect 385 138 401 172
rect 489 138 505 172
rect 563 138 579 172
rect 667 138 683 172
rect 741 138 757 172
rect 845 138 861 172
rect -907 88 -873 104
rect -907 -104 -873 -88
rect -729 88 -695 104
rect -729 -104 -695 -88
rect -551 88 -517 104
rect -551 -104 -517 -88
rect -373 88 -339 104
rect -373 -104 -339 -88
rect -195 88 -161 104
rect -195 -104 -161 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 161 88 195 104
rect 161 -104 195 -88
rect 339 88 373 104
rect 339 -104 373 -88
rect 517 88 551 104
rect 517 -104 551 -88
rect 695 88 729 104
rect 695 -104 729 -88
rect 873 88 907 104
rect 873 -104 907 -88
rect -861 -172 -845 -138
rect -757 -172 -741 -138
rect -683 -172 -667 -138
rect -579 -172 -563 -138
rect -505 -172 -489 -138
rect -401 -172 -385 -138
rect -327 -172 -311 -138
rect -223 -172 -207 -138
rect -149 -172 -133 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 133 -172 149 -138
rect 207 -172 223 -138
rect 311 -172 327 -138
rect 385 -172 401 -138
rect 489 -172 505 -138
rect 563 -172 579 -138
rect 667 -172 683 -138
rect 741 -172 757 -138
rect 845 -172 861 -138
rect -1021 -240 -987 -178
rect 987 -240 1021 -178
rect -1021 -274 -925 -240
rect 925 -274 1021 -240
<< viali >>
rect -845 138 -757 172
rect -667 138 -579 172
rect -489 138 -401 172
rect -311 138 -223 172
rect -133 138 -45 172
rect 45 138 133 172
rect 223 138 311 172
rect 401 138 489 172
rect 579 138 667 172
rect 757 138 845 172
rect -907 -88 -873 88
rect -729 -88 -695 88
rect -551 -88 -517 88
rect -373 -88 -339 88
rect -195 -88 -161 88
rect -17 -88 17 88
rect 161 -88 195 88
rect 339 -88 373 88
rect 517 -88 551 88
rect 695 -88 729 88
rect 873 -88 907 88
rect -845 -172 -757 -138
rect -667 -172 -579 -138
rect -489 -172 -401 -138
rect -311 -172 -223 -138
rect -133 -172 -45 -138
rect 45 -172 133 -138
rect 223 -172 311 -138
rect 401 -172 489 -138
rect 579 -172 667 -138
rect 757 -172 845 -138
<< metal1 >>
rect -857 172 -745 178
rect -857 138 -845 172
rect -757 138 -745 172
rect -857 132 -745 138
rect -679 172 -567 178
rect -679 138 -667 172
rect -579 138 -567 172
rect -679 132 -567 138
rect -501 172 -389 178
rect -501 138 -489 172
rect -401 138 -389 172
rect -501 132 -389 138
rect -323 172 -211 178
rect -323 138 -311 172
rect -223 138 -211 172
rect -323 132 -211 138
rect -145 172 -33 178
rect -145 138 -133 172
rect -45 138 -33 172
rect -145 132 -33 138
rect 33 172 145 178
rect 33 138 45 172
rect 133 138 145 172
rect 33 132 145 138
rect 211 172 323 178
rect 211 138 223 172
rect 311 138 323 172
rect 211 132 323 138
rect 389 172 501 178
rect 389 138 401 172
rect 489 138 501 172
rect 389 132 501 138
rect 567 172 679 178
rect 567 138 579 172
rect 667 138 679 172
rect 567 132 679 138
rect 745 172 857 178
rect 745 138 757 172
rect 845 138 857 172
rect 745 132 857 138
rect -913 88 -867 100
rect -913 -88 -907 88
rect -873 -88 -867 88
rect -913 -100 -867 -88
rect -735 88 -689 100
rect -735 -88 -729 88
rect -695 -88 -689 88
rect -735 -100 -689 -88
rect -557 88 -511 100
rect -557 -88 -551 88
rect -517 -88 -511 88
rect -557 -100 -511 -88
rect -379 88 -333 100
rect -379 -88 -373 88
rect -339 -88 -333 88
rect -379 -100 -333 -88
rect -201 88 -155 100
rect -201 -88 -195 88
rect -161 -88 -155 88
rect -201 -100 -155 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 155 88 201 100
rect 155 -88 161 88
rect 195 -88 201 88
rect 155 -100 201 -88
rect 333 88 379 100
rect 333 -88 339 88
rect 373 -88 379 88
rect 333 -100 379 -88
rect 511 88 557 100
rect 511 -88 517 88
rect 551 -88 557 88
rect 511 -100 557 -88
rect 689 88 735 100
rect 689 -88 695 88
rect 729 -88 735 88
rect 689 -100 735 -88
rect 867 88 913 100
rect 867 -88 873 88
rect 907 -88 913 88
rect 867 -100 913 -88
rect -857 -138 -745 -132
rect -857 -172 -845 -138
rect -757 -172 -745 -138
rect -857 -178 -745 -172
rect -679 -138 -567 -132
rect -679 -172 -667 -138
rect -579 -172 -567 -138
rect -679 -178 -567 -172
rect -501 -138 -389 -132
rect -501 -172 -489 -138
rect -401 -172 -389 -138
rect -501 -178 -389 -172
rect -323 -138 -211 -132
rect -323 -172 -311 -138
rect -223 -172 -211 -138
rect -323 -178 -211 -172
rect -145 -138 -33 -132
rect -145 -172 -133 -138
rect -45 -172 -33 -138
rect -145 -178 -33 -172
rect 33 -138 145 -132
rect 33 -172 45 -138
rect 133 -172 145 -138
rect 33 -178 145 -172
rect 211 -138 323 -132
rect 211 -172 223 -138
rect 311 -172 323 -138
rect 211 -178 323 -172
rect 389 -138 501 -132
rect 389 -172 401 -138
rect 489 -172 501 -138
rect 389 -178 501 -172
rect 567 -138 679 -132
rect 567 -172 579 -138
rect 667 -172 679 -138
rect 567 -178 679 -172
rect 745 -138 857 -132
rect 745 -172 757 -138
rect 845 -172 857 -138
rect 745 -178 857 -172
<< properties >>
string FIXED_BBOX -1004 -257 1004 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.6 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
