magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -365 162 -307 168
rect -173 162 -115 168
rect 19 162 77 168
rect 211 162 269 168
rect 403 162 461 168
rect -365 128 -353 162
rect -173 128 -161 162
rect 19 128 31 162
rect 211 128 223 162
rect 403 128 415 162
rect -365 122 -307 128
rect -173 122 -115 128
rect 19 122 77 128
rect 211 122 269 128
rect 403 122 461 128
rect -461 -128 -403 -122
rect -269 -128 -211 -122
rect -77 -128 -19 -122
rect 115 -128 173 -122
rect 307 -128 365 -122
rect -461 -162 -449 -128
rect -269 -162 -257 -128
rect -77 -162 -65 -128
rect 115 -162 127 -128
rect 307 -162 319 -128
rect -461 -168 -403 -162
rect -269 -168 -211 -162
rect -77 -168 -19 -162
rect 115 -168 173 -162
rect 307 -168 365 -162
<< pwell >>
rect -647 -300 647 300
<< nmos >>
rect -447 -90 -417 90
rect -351 -90 -321 90
rect -255 -90 -225 90
rect -159 -90 -129 90
rect -63 -90 -33 90
rect 33 -90 63 90
rect 129 -90 159 90
rect 225 -90 255 90
rect 321 -90 351 90
rect 417 -90 447 90
<< ndiff >>
rect -509 78 -447 90
rect -509 -78 -497 78
rect -463 -78 -447 78
rect -509 -90 -447 -78
rect -417 78 -351 90
rect -417 -78 -401 78
rect -367 -78 -351 78
rect -417 -90 -351 -78
rect -321 78 -255 90
rect -321 -78 -305 78
rect -271 -78 -255 78
rect -321 -90 -255 -78
rect -225 78 -159 90
rect -225 -78 -209 78
rect -175 -78 -159 78
rect -225 -90 -159 -78
rect -129 78 -63 90
rect -129 -78 -113 78
rect -79 -78 -63 78
rect -129 -90 -63 -78
rect -33 78 33 90
rect -33 -78 -17 78
rect 17 -78 33 78
rect -33 -90 33 -78
rect 63 78 129 90
rect 63 -78 79 78
rect 113 -78 129 78
rect 63 -90 129 -78
rect 159 78 225 90
rect 159 -78 175 78
rect 209 -78 225 78
rect 159 -90 225 -78
rect 255 78 321 90
rect 255 -78 271 78
rect 305 -78 321 78
rect 255 -90 321 -78
rect 351 78 417 90
rect 351 -78 367 78
rect 401 -78 417 78
rect 351 -90 417 -78
rect 447 78 509 90
rect 447 -78 463 78
rect 497 -78 509 78
rect 447 -90 509 -78
<< ndiffc >>
rect -497 -78 -463 78
rect -401 -78 -367 78
rect -305 -78 -271 78
rect -209 -78 -175 78
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
rect 175 -78 209 78
rect 271 -78 305 78
rect 367 -78 401 78
rect 463 -78 497 78
<< psubdiff >>
rect -611 230 -515 264
rect 515 230 611 264
rect -611 168 -577 230
rect 577 168 611 230
rect -611 -230 -577 -168
rect 577 -230 611 -168
rect -611 -264 -515 -230
rect 515 -264 611 -230
<< psubdiffcont >>
rect -515 230 515 264
rect -611 -168 -577 168
rect 577 -168 611 168
rect -515 -264 515 -230
<< poly >>
rect -369 162 -303 178
rect -369 128 -353 162
rect -319 128 -303 162
rect -447 90 -417 116
rect -369 112 -303 128
rect -177 162 -111 178
rect -177 128 -161 162
rect -127 128 -111 162
rect -351 90 -321 112
rect -255 90 -225 116
rect -177 112 -111 128
rect 15 162 81 178
rect 15 128 31 162
rect 65 128 81 162
rect -159 90 -129 112
rect -63 90 -33 116
rect 15 112 81 128
rect 207 162 273 178
rect 207 128 223 162
rect 257 128 273 162
rect 33 90 63 112
rect 129 90 159 116
rect 207 112 273 128
rect 399 162 465 178
rect 399 128 415 162
rect 449 128 465 162
rect 225 90 255 112
rect 321 90 351 116
rect 399 112 465 128
rect 417 90 447 112
rect -447 -112 -417 -90
rect -465 -128 -399 -112
rect -351 -116 -321 -90
rect -255 -112 -225 -90
rect -465 -162 -449 -128
rect -415 -162 -399 -128
rect -465 -178 -399 -162
rect -273 -128 -207 -112
rect -159 -116 -129 -90
rect -63 -112 -33 -90
rect -273 -162 -257 -128
rect -223 -162 -207 -128
rect -273 -178 -207 -162
rect -81 -128 -15 -112
rect 33 -116 63 -90
rect 129 -112 159 -90
rect -81 -162 -65 -128
rect -31 -162 -15 -128
rect -81 -178 -15 -162
rect 111 -128 177 -112
rect 225 -116 255 -90
rect 321 -112 351 -90
rect 111 -162 127 -128
rect 161 -162 177 -128
rect 111 -178 177 -162
rect 303 -128 369 -112
rect 417 -116 447 -90
rect 303 -162 319 -128
rect 353 -162 369 -128
rect 303 -178 369 -162
<< polycont >>
rect -353 128 -319 162
rect -161 128 -127 162
rect 31 128 65 162
rect 223 128 257 162
rect 415 128 449 162
rect -449 -162 -415 -128
rect -257 -162 -223 -128
rect -65 -162 -31 -128
rect 127 -162 161 -128
rect 319 -162 353 -128
<< locali >>
rect -611 230 -515 264
rect 515 230 611 264
rect -611 168 -577 230
rect 577 168 611 230
rect -369 128 -353 162
rect -319 128 -303 162
rect -177 128 -161 162
rect -127 128 -111 162
rect 15 128 31 162
rect 65 128 81 162
rect 207 128 223 162
rect 257 128 273 162
rect 399 128 415 162
rect 449 128 465 162
rect -497 78 -463 94
rect -497 -94 -463 -78
rect -401 78 -367 94
rect -401 -94 -367 -78
rect -305 78 -271 94
rect -305 -94 -271 -78
rect -209 78 -175 94
rect -209 -94 -175 -78
rect -113 78 -79 94
rect -113 -94 -79 -78
rect -17 78 17 94
rect -17 -94 17 -78
rect 79 78 113 94
rect 79 -94 113 -78
rect 175 78 209 94
rect 175 -94 209 -78
rect 271 78 305 94
rect 271 -94 305 -78
rect 367 78 401 94
rect 367 -94 401 -78
rect 463 78 497 94
rect 463 -94 497 -78
rect -465 -162 -449 -128
rect -415 -162 -399 -128
rect -273 -162 -257 -128
rect -223 -162 -207 -128
rect -81 -162 -65 -128
rect -31 -162 -15 -128
rect 111 -162 127 -128
rect 161 -162 177 -128
rect 303 -162 319 -128
rect 353 -162 369 -128
rect -611 -230 -577 -168
rect 577 -230 611 -168
rect -611 -264 -515 -230
rect 515 -264 611 -230
<< viali >>
rect -353 128 -319 162
rect -161 128 -127 162
rect 31 128 65 162
rect 223 128 257 162
rect 415 128 449 162
rect -497 -78 -463 78
rect -401 -78 -367 78
rect -305 -78 -271 78
rect -209 -78 -175 78
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
rect 175 -78 209 78
rect 271 -78 305 78
rect 367 -78 401 78
rect 463 -78 497 78
rect -449 -162 -415 -128
rect -257 -162 -223 -128
rect -65 -162 -31 -128
rect 127 -162 161 -128
rect 319 -162 353 -128
<< metal1 >>
rect -365 162 -307 168
rect -365 128 -353 162
rect -319 128 -307 162
rect -365 122 -307 128
rect -173 162 -115 168
rect -173 128 -161 162
rect -127 128 -115 162
rect -173 122 -115 128
rect 19 162 77 168
rect 19 128 31 162
rect 65 128 77 162
rect 19 122 77 128
rect 211 162 269 168
rect 211 128 223 162
rect 257 128 269 162
rect 211 122 269 128
rect 403 162 461 168
rect 403 128 415 162
rect 449 128 461 162
rect 403 122 461 128
rect -503 78 -457 90
rect -503 -78 -497 78
rect -463 -78 -457 78
rect -503 -90 -457 -78
rect -407 78 -361 90
rect -407 -78 -401 78
rect -367 -78 -361 78
rect -407 -90 -361 -78
rect -311 78 -265 90
rect -311 -78 -305 78
rect -271 -78 -265 78
rect -311 -90 -265 -78
rect -215 78 -169 90
rect -215 -78 -209 78
rect -175 -78 -169 78
rect -215 -90 -169 -78
rect -119 78 -73 90
rect -119 -78 -113 78
rect -79 -78 -73 78
rect -119 -90 -73 -78
rect -23 78 23 90
rect -23 -78 -17 78
rect 17 -78 23 78
rect -23 -90 23 -78
rect 73 78 119 90
rect 73 -78 79 78
rect 113 -78 119 78
rect 73 -90 119 -78
rect 169 78 215 90
rect 169 -78 175 78
rect 209 -78 215 78
rect 169 -90 215 -78
rect 265 78 311 90
rect 265 -78 271 78
rect 305 -78 311 78
rect 265 -90 311 -78
rect 361 78 407 90
rect 361 -78 367 78
rect 401 -78 407 78
rect 361 -90 407 -78
rect 457 78 503 90
rect 457 -78 463 78
rect 497 -78 503 78
rect 457 -90 503 -78
rect -461 -128 -403 -122
rect -461 -162 -449 -128
rect -415 -162 -403 -128
rect -461 -168 -403 -162
rect -269 -128 -211 -122
rect -269 -162 -257 -128
rect -223 -162 -211 -128
rect -269 -168 -211 -162
rect -77 -128 -19 -122
rect -77 -162 -65 -128
rect -31 -162 -19 -128
rect -77 -168 -19 -162
rect 115 -128 173 -122
rect 115 -162 127 -128
rect 161 -162 173 -128
rect 115 -168 173 -162
rect 307 -128 365 -122
rect 307 -162 319 -128
rect 353 -162 365 -128
rect 307 -168 365 -162
<< properties >>
string FIXED_BBOX -594 -247 594 247
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.9 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
