magic
tech sky130A
magscale 1 2
timestamp 1707817411
<< error_p >>
rect -29 681 29 687
rect -29 647 -17 681
rect -29 641 29 647
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect -29 -687 29 -681
<< nwell >>
rect -226 -819 226 819
<< pmos >>
rect -30 -600 30 600
<< pdiff >>
rect -88 588 -30 600
rect -88 -588 -76 588
rect -42 -588 -30 588
rect -88 -600 -30 -588
rect 30 588 88 600
rect 30 -588 42 588
rect 76 -588 88 588
rect 30 -600 88 -588
<< pdiffc >>
rect -76 -588 -42 588
rect 42 -588 76 588
<< nsubdiff >>
rect -190 749 -94 783
rect 94 749 190 783
rect -190 687 -156 749
rect 156 687 190 749
rect -190 -749 -156 -687
rect 156 -749 190 -687
rect -190 -783 -94 -749
rect 94 -783 190 -749
<< nsubdiffcont >>
rect -94 749 94 783
rect -190 -687 -156 687
rect 156 -687 190 687
rect -94 -783 94 -749
<< poly >>
rect -33 681 33 697
rect -33 647 -17 681
rect 17 647 33 681
rect -33 631 33 647
rect -30 600 30 631
rect -30 -631 30 -600
rect -33 -647 33 -631
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -697 33 -681
<< polycont >>
rect -17 647 17 681
rect -17 -681 17 -647
<< locali >>
rect -190 749 -94 783
rect 94 749 190 783
rect -190 687 -156 749
rect 156 687 190 749
rect -33 647 -17 681
rect 17 647 33 681
rect -76 588 -42 604
rect -76 -604 -42 -588
rect 42 588 76 604
rect 42 -604 76 -588
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -190 -749 -156 -687
rect 156 -749 190 -687
rect -190 -783 -94 -749
rect 94 -783 190 -749
<< viali >>
rect -17 647 17 681
rect -76 -588 -42 588
rect 42 -588 76 588
rect -17 -681 17 -647
<< metal1 >>
rect -29 681 29 687
rect -29 647 -17 681
rect 17 647 29 681
rect -29 641 29 647
rect -82 588 -36 600
rect -82 -588 -76 588
rect -42 -588 -36 588
rect -82 -600 -36 -588
rect 36 588 82 600
rect 36 -588 42 588
rect 76 -588 82 588
rect 36 -600 82 -588
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect 17 -681 29 -647
rect -29 -687 29 -681
<< properties >>
string FIXED_BBOX -173 -766 173 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
