magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -125 672 -67 678
rect 67 672 125 678
rect -125 638 -113 672
rect 67 638 79 672
rect -125 632 -67 638
rect 67 632 125 638
rect -221 -638 -163 -632
rect -29 -638 29 -632
rect 163 -638 221 -632
rect -221 -672 -209 -638
rect -29 -672 -17 -638
rect 163 -672 175 -638
rect -221 -678 -163 -672
rect -29 -678 29 -672
rect 163 -678 221 -672
<< pwell >>
rect -407 -810 407 810
<< nmos >>
rect -207 -600 -177 600
rect -111 -600 -81 600
rect -15 -600 15 600
rect 81 -600 111 600
rect 177 -600 207 600
<< ndiff >>
rect -269 588 -207 600
rect -269 -588 -257 588
rect -223 -588 -207 588
rect -269 -600 -207 -588
rect -177 588 -111 600
rect -177 -588 -161 588
rect -127 -588 -111 588
rect -177 -600 -111 -588
rect -81 588 -15 600
rect -81 -588 -65 588
rect -31 -588 -15 588
rect -81 -600 -15 -588
rect 15 588 81 600
rect 15 -588 31 588
rect 65 -588 81 588
rect 15 -600 81 -588
rect 111 588 177 600
rect 111 -588 127 588
rect 161 -588 177 588
rect 111 -600 177 -588
rect 207 588 269 600
rect 207 -588 223 588
rect 257 -588 269 588
rect 207 -600 269 -588
<< ndiffc >>
rect -257 -588 -223 588
rect -161 -588 -127 588
rect -65 -588 -31 588
rect 31 -588 65 588
rect 127 -588 161 588
rect 223 -588 257 588
<< psubdiff >>
rect -371 740 -275 774
rect 275 740 371 774
rect -371 678 -337 740
rect 337 678 371 740
rect -371 -740 -337 -678
rect 337 -740 371 -678
rect -371 -774 -275 -740
rect 275 -774 371 -740
<< psubdiffcont >>
rect -275 740 275 774
rect -371 -678 -337 678
rect 337 -678 371 678
rect -275 -774 275 -740
<< poly >>
rect -129 672 -63 688
rect -129 638 -113 672
rect -79 638 -63 672
rect -207 600 -177 626
rect -129 622 -63 638
rect 63 672 129 688
rect 63 638 79 672
rect 113 638 129 672
rect -111 600 -81 622
rect -15 600 15 626
rect 63 622 129 638
rect 81 600 111 622
rect 177 600 207 626
rect -207 -622 -177 -600
rect -225 -638 -159 -622
rect -111 -626 -81 -600
rect -15 -622 15 -600
rect -225 -672 -209 -638
rect -175 -672 -159 -638
rect -225 -688 -159 -672
rect -33 -638 33 -622
rect 81 -626 111 -600
rect 177 -622 207 -600
rect -33 -672 -17 -638
rect 17 -672 33 -638
rect -33 -688 33 -672
rect 159 -638 225 -622
rect 159 -672 175 -638
rect 209 -672 225 -638
rect 159 -688 225 -672
<< polycont >>
rect -113 638 -79 672
rect 79 638 113 672
rect -209 -672 -175 -638
rect -17 -672 17 -638
rect 175 -672 209 -638
<< locali >>
rect -371 740 -275 774
rect 275 740 371 774
rect -371 678 -337 740
rect 337 678 371 740
rect -129 638 -113 672
rect -79 638 -63 672
rect 63 638 79 672
rect 113 638 129 672
rect -257 588 -223 604
rect -257 -604 -223 -588
rect -161 588 -127 604
rect -161 -604 -127 -588
rect -65 588 -31 604
rect -65 -604 -31 -588
rect 31 588 65 604
rect 31 -604 65 -588
rect 127 588 161 604
rect 127 -604 161 -588
rect 223 588 257 604
rect 223 -604 257 -588
rect -225 -672 -209 -638
rect -175 -672 -159 -638
rect -33 -672 -17 -638
rect 17 -672 33 -638
rect 159 -672 175 -638
rect 209 -672 225 -638
rect -371 -740 -337 -678
rect 337 -740 371 -678
rect -371 -774 -275 -740
rect 275 -774 371 -740
<< viali >>
rect -113 638 -79 672
rect 79 638 113 672
rect -257 -588 -223 588
rect -161 -588 -127 588
rect -65 -588 -31 588
rect 31 -588 65 588
rect 127 -588 161 588
rect 223 -588 257 588
rect -209 -672 -175 -638
rect -17 -672 17 -638
rect 175 -672 209 -638
<< metal1 >>
rect -125 672 -67 678
rect -125 638 -113 672
rect -79 638 -67 672
rect -125 632 -67 638
rect 67 672 125 678
rect 67 638 79 672
rect 113 638 125 672
rect 67 632 125 638
rect -263 588 -217 600
rect -263 -588 -257 588
rect -223 -588 -217 588
rect -263 -600 -217 -588
rect -167 588 -121 600
rect -167 -588 -161 588
rect -127 -588 -121 588
rect -167 -600 -121 -588
rect -71 588 -25 600
rect -71 -588 -65 588
rect -31 -588 -25 588
rect -71 -600 -25 -588
rect 25 588 71 600
rect 25 -588 31 588
rect 65 -588 71 588
rect 25 -600 71 -588
rect 121 588 167 600
rect 121 -588 127 588
rect 161 -588 167 588
rect 121 -600 167 -588
rect 217 588 263 600
rect 217 -588 223 588
rect 257 -588 263 588
rect 217 -600 263 -588
rect -221 -638 -163 -632
rect -221 -672 -209 -638
rect -175 -672 -163 -638
rect -221 -678 -163 -672
rect -29 -638 29 -632
rect -29 -672 -17 -638
rect 17 -672 29 -638
rect -29 -678 29 -672
rect 163 -638 221 -632
rect 163 -672 175 -638
rect 209 -672 221 -638
rect 163 -678 221 -672
<< properties >>
string FIXED_BBOX -354 -757 354 757
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
