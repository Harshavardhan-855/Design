magic
tech sky130A
magscale 1 2
timestamp 1709102441
<< error_p >>
rect -365 981 -307 987
rect -173 981 -115 987
rect 19 981 77 987
rect 211 981 269 987
rect 403 981 461 987
rect -365 947 -353 981
rect -173 947 -161 981
rect 19 947 31 981
rect 211 947 223 981
rect 403 947 415 981
rect -365 941 -307 947
rect -173 941 -115 947
rect 19 941 77 947
rect 211 941 269 947
rect 403 941 461 947
rect -461 -947 -403 -941
rect -269 -947 -211 -941
rect -77 -947 -19 -941
rect 115 -947 173 -941
rect 307 -947 365 -941
rect -461 -981 -449 -947
rect -269 -981 -257 -947
rect -77 -981 -65 -947
rect 115 -981 127 -947
rect 307 -981 319 -947
rect -461 -987 -403 -981
rect -269 -987 -211 -981
rect -77 -987 -19 -981
rect 115 -987 173 -981
rect 307 -987 365 -981
<< nwell >>
rect -647 -1119 647 1119
<< pmos >>
rect -447 -900 -417 900
rect -351 -900 -321 900
rect -255 -900 -225 900
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
rect 225 -900 255 900
rect 321 -900 351 900
rect 417 -900 447 900
<< pdiff >>
rect -509 888 -447 900
rect -509 -888 -497 888
rect -463 -888 -447 888
rect -509 -900 -447 -888
rect -417 888 -351 900
rect -417 -888 -401 888
rect -367 -888 -351 888
rect -417 -900 -351 -888
rect -321 888 -255 900
rect -321 -888 -305 888
rect -271 -888 -255 888
rect -321 -900 -255 -888
rect -225 888 -159 900
rect -225 -888 -209 888
rect -175 -888 -159 888
rect -225 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 225 900
rect 159 -888 175 888
rect 209 -888 225 888
rect 159 -900 225 -888
rect 255 888 321 900
rect 255 -888 271 888
rect 305 -888 321 888
rect 255 -900 321 -888
rect 351 888 417 900
rect 351 -888 367 888
rect 401 -888 417 888
rect 351 -900 417 -888
rect 447 888 509 900
rect 447 -888 463 888
rect 497 -888 509 888
rect 447 -900 509 -888
<< pdiffc >>
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
<< nsubdiff >>
rect -611 1049 -515 1083
rect 515 1049 611 1083
rect -611 987 -577 1049
rect 577 987 611 1049
rect -611 -1049 -577 -987
rect 577 -1049 611 -987
rect -611 -1083 -515 -1049
rect 515 -1083 611 -1049
<< nsubdiffcont >>
rect -515 1049 515 1083
rect -611 -987 -577 987
rect 577 -987 611 987
rect -515 -1083 515 -1049
<< poly >>
rect -369 981 -303 997
rect -369 947 -353 981
rect -319 947 -303 981
rect -369 931 -303 947
rect -177 981 -111 997
rect -177 947 -161 981
rect -127 947 -111 981
rect -177 931 -111 947
rect 15 981 81 997
rect 15 947 31 981
rect 65 947 81 981
rect 15 931 81 947
rect 207 981 273 997
rect 207 947 223 981
rect 257 947 273 981
rect 207 931 273 947
rect 399 981 465 997
rect 399 947 415 981
rect 449 947 465 981
rect 399 931 465 947
rect -447 900 -417 926
rect -351 900 -321 931
rect -255 900 -225 926
rect -159 900 -129 931
rect -63 900 -33 926
rect 33 900 63 931
rect 129 900 159 926
rect 225 900 255 931
rect 321 900 351 926
rect 417 900 447 931
rect -447 -931 -417 -900
rect -351 -926 -321 -900
rect -255 -931 -225 -900
rect -159 -926 -129 -900
rect -63 -931 -33 -900
rect 33 -926 63 -900
rect 129 -931 159 -900
rect 225 -926 255 -900
rect 321 -931 351 -900
rect 417 -926 447 -900
rect -465 -947 -399 -931
rect -465 -981 -449 -947
rect -415 -981 -399 -947
rect -465 -997 -399 -981
rect -273 -947 -207 -931
rect -273 -981 -257 -947
rect -223 -981 -207 -947
rect -273 -997 -207 -981
rect -81 -947 -15 -931
rect -81 -981 -65 -947
rect -31 -981 -15 -947
rect -81 -997 -15 -981
rect 111 -947 177 -931
rect 111 -981 127 -947
rect 161 -981 177 -947
rect 111 -997 177 -981
rect 303 -947 369 -931
rect 303 -981 319 -947
rect 353 -981 369 -947
rect 303 -997 369 -981
<< polycont >>
rect -353 947 -319 981
rect -161 947 -127 981
rect 31 947 65 981
rect 223 947 257 981
rect 415 947 449 981
rect -449 -981 -415 -947
rect -257 -981 -223 -947
rect -65 -981 -31 -947
rect 127 -981 161 -947
rect 319 -981 353 -947
<< locali >>
rect -611 1049 -515 1083
rect 515 1049 611 1083
rect -611 987 -577 1049
rect 577 987 611 1049
rect -369 947 -353 981
rect -319 947 -303 981
rect -177 947 -161 981
rect -127 947 -111 981
rect 15 947 31 981
rect 65 947 81 981
rect 207 947 223 981
rect 257 947 273 981
rect 399 947 415 981
rect 449 947 465 981
rect -497 888 -463 904
rect -497 -904 -463 -888
rect -401 888 -367 904
rect -401 -904 -367 -888
rect -305 888 -271 904
rect -305 -904 -271 -888
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect 271 888 305 904
rect 271 -904 305 -888
rect 367 888 401 904
rect 367 -904 401 -888
rect 463 888 497 904
rect 463 -904 497 -888
rect -465 -981 -449 -947
rect -415 -981 -399 -947
rect -273 -981 -257 -947
rect -223 -981 -207 -947
rect -81 -981 -65 -947
rect -31 -981 -15 -947
rect 111 -981 127 -947
rect 161 -981 177 -947
rect 303 -981 319 -947
rect 353 -981 369 -947
rect -611 -1049 -577 -987
rect 577 -1049 611 -987
rect -611 -1083 -515 -1049
rect 515 -1083 611 -1049
<< viali >>
rect -353 947 -319 981
rect -161 947 -127 981
rect 31 947 65 981
rect 223 947 257 981
rect 415 947 449 981
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect -449 -981 -415 -947
rect -257 -981 -223 -947
rect -65 -981 -31 -947
rect 127 -981 161 -947
rect 319 -981 353 -947
<< metal1 >>
rect -365 981 -307 987
rect -365 947 -353 981
rect -319 947 -307 981
rect -365 941 -307 947
rect -173 981 -115 987
rect -173 947 -161 981
rect -127 947 -115 981
rect -173 941 -115 947
rect 19 981 77 987
rect 19 947 31 981
rect 65 947 77 981
rect 19 941 77 947
rect 211 981 269 987
rect 211 947 223 981
rect 257 947 269 981
rect 211 941 269 947
rect 403 981 461 987
rect 403 947 415 981
rect 449 947 461 981
rect 403 941 461 947
rect -503 888 -457 900
rect -503 -888 -497 888
rect -463 -888 -457 888
rect -503 -900 -457 -888
rect -407 888 -361 900
rect -407 -888 -401 888
rect -367 -888 -361 888
rect -407 -900 -361 -888
rect -311 888 -265 900
rect -311 -888 -305 888
rect -271 -888 -265 888
rect -311 -900 -265 -888
rect -215 888 -169 900
rect -215 -888 -209 888
rect -175 -888 -169 888
rect -215 -900 -169 -888
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 169 888 215 900
rect 169 -888 175 888
rect 209 -888 215 888
rect 169 -900 215 -888
rect 265 888 311 900
rect 265 -888 271 888
rect 305 -888 311 888
rect 265 -900 311 -888
rect 361 888 407 900
rect 361 -888 367 888
rect 401 -888 407 888
rect 361 -900 407 -888
rect 457 888 503 900
rect 457 -888 463 888
rect 497 -888 503 888
rect 457 -900 503 -888
rect -461 -947 -403 -941
rect -461 -981 -449 -947
rect -415 -981 -403 -947
rect -461 -987 -403 -981
rect -269 -947 -211 -941
rect -269 -981 -257 -947
rect -223 -981 -211 -947
rect -269 -987 -211 -981
rect -77 -947 -19 -941
rect -77 -981 -65 -947
rect -31 -981 -19 -947
rect -77 -987 -19 -981
rect 115 -947 173 -941
rect 115 -981 127 -947
rect 161 -981 173 -947
rect 115 -987 173 -981
rect 307 -947 365 -941
rect 307 -981 319 -947
rect 353 -981 365 -947
rect 307 -987 365 -981
<< properties >>
string FIXED_BBOX -594 -1066 594 1066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
