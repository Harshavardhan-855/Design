magic
tech sky130A
magscale 1 2
timestamp 1706848405
<< viali >>
rect 2710 1624 2840 1672
rect 3652 1626 3796 1688
rect 4844 892 4968 1056
rect 5338 490 5484 582
rect 2234 -1228 2332 -1176
rect 3992 -1224 4112 -1178
rect 2264 -1650 2342 -1572
rect 3974 -1648 4178 -1578
rect 3088 -2760 3526 -2596
<< metal1 >>
rect 3210 1952 3410 2008
rect 3210 1866 3270 1952
rect 3352 1866 3410 1952
rect 3210 1808 3410 1866
rect 2668 1610 2678 1684
rect 2864 1610 2874 1684
rect 3614 1616 3624 1708
rect 3820 1616 3830 1708
rect 1852 1566 2996 1574
rect 3622 1566 4766 1580
rect 1852 1520 4766 1566
rect 1852 1514 2996 1520
rect 1806 1244 1816 1448
rect 1876 1244 1886 1448
rect 2042 1252 2052 1456
rect 2112 1252 2122 1456
rect 2276 1248 2286 1452
rect 2346 1248 2356 1452
rect 2514 1252 2524 1456
rect 2584 1252 2594 1456
rect 2750 1260 2760 1464
rect 2820 1260 2830 1464
rect 2988 1266 2998 1470
rect 3058 1266 3068 1470
rect 1908 506 1918 710
rect 1978 506 1988 710
rect 2144 512 2154 716
rect 2214 512 2224 716
rect 2382 512 2392 716
rect 2452 512 2462 716
rect 2620 512 2630 716
rect 2690 512 2700 716
rect 3276 712 3342 1520
rect 3558 1222 3568 1444
rect 3630 1222 3640 1444
rect 3794 1216 3804 1438
rect 3866 1216 3876 1438
rect 4032 1220 4042 1442
rect 4104 1220 4114 1442
rect 4266 1224 4276 1446
rect 4338 1224 4348 1446
rect 4500 1224 4510 1446
rect 4572 1224 4582 1446
rect 4742 1234 4752 1456
rect 4814 1234 4824 1456
rect 4838 1056 4974 1068
rect 4838 892 4844 1056
rect 4968 1022 4974 1056
rect 4968 1018 5442 1022
rect 4968 912 5450 1018
rect 4968 892 4974 912
rect 4838 880 4974 892
rect 2854 508 2864 712
rect 2924 508 2934 712
rect 3270 526 3280 712
rect 3338 526 3348 712
rect 1854 430 2998 444
rect 3276 430 3342 526
rect 3684 498 3694 720
rect 3756 498 3766 720
rect 3922 504 3932 726
rect 3994 504 4004 726
rect 4156 508 4166 730
rect 4228 508 4238 730
rect 4388 510 4398 732
rect 4460 510 4470 732
rect 4632 598 4642 732
rect 4630 510 4642 598
rect 4704 598 4714 732
rect 5336 610 5450 912
rect 4704 510 4722 598
rect 5280 488 5290 610
rect 5520 488 5530 610
rect 5326 484 5496 488
rect 3622 444 4630 446
rect 4722 444 4766 446
rect 3622 430 4766 444
rect 1854 394 4766 430
rect 5096 398 6552 456
rect 1854 386 4630 394
rect 4722 386 4766 394
rect 1854 384 3708 386
rect 3276 382 3342 384
rect 5098 272 5182 398
rect 5408 396 6552 398
rect 5090 126 5100 272
rect 5178 126 5188 272
rect 3622 60 4630 62
rect 4722 60 4766 62
rect 3622 52 4766 60
rect 1852 42 2996 44
rect 1404 -10 2996 42
rect 3324 2 4766 52
rect 3324 -2 3680 2
rect 4624 0 4762 2
rect 1450 -468 1506 -10
rect 1852 -16 2996 -10
rect 1794 -308 1804 -74
rect 1868 -308 1878 -74
rect 2032 -304 2042 -70
rect 2106 -304 2116 -70
rect 2266 -296 2276 -62
rect 2340 -296 2350 -62
rect 2504 -292 2514 -58
rect 2578 -292 2588 -58
rect 2738 -290 2748 -56
rect 2812 -290 2822 -56
rect 2976 -290 2986 -56
rect 3050 -290 3060 -56
rect 1288 -668 1506 -468
rect 1450 -1082 1506 -668
rect 1914 -1034 1924 -800
rect 1988 -1034 1998 -800
rect 2148 -1034 2158 -800
rect 2222 -1034 2232 -800
rect 2388 -1032 2398 -798
rect 2462 -1032 2472 -798
rect 2622 -1032 2632 -798
rect 2696 -1032 2706 -798
rect 2860 -1028 2870 -794
rect 2934 -1028 2944 -794
rect 3326 -1054 3386 -2
rect 3568 -362 3578 -108
rect 3630 -362 3640 -108
rect 3798 -362 3808 -114
rect 3864 -362 3874 -114
rect 4034 -356 4044 -108
rect 4100 -356 4110 -108
rect 4274 -348 4284 -100
rect 4340 -348 4350 -100
rect 4510 -336 4520 -88
rect 4576 -336 4586 -88
rect 4744 -330 4754 -82
rect 4810 -330 4820 -82
rect 5098 -680 5182 126
rect 5354 100 5364 310
rect 5432 100 5442 310
rect 5592 100 5602 310
rect 5670 100 5680 310
rect 5836 104 5846 314
rect 5914 104 5924 314
rect 6066 104 6076 314
rect 6144 104 6154 314
rect 6304 108 6314 318
rect 6382 108 6392 318
rect 6536 106 6546 316
rect 6614 106 6624 316
rect 5474 -622 5484 -412
rect 5552 -622 5562 -412
rect 5708 -618 5718 -408
rect 5786 -618 5796 -408
rect 5946 -620 5956 -410
rect 6024 -620 6034 -410
rect 6178 -624 6188 -414
rect 6256 -624 6266 -414
rect 6418 -618 6428 -408
rect 6496 -618 6506 -408
rect 5364 -680 6508 -678
rect 5098 -738 6508 -680
rect 5098 -740 5400 -738
rect 3684 -1002 3694 -774
rect 3760 -1002 3770 -774
rect 3922 -1000 3932 -772
rect 3998 -1000 4008 -772
rect 4160 -1002 4170 -774
rect 4236 -1002 4246 -774
rect 4398 -1002 4408 -774
rect 4474 -1002 4484 -774
rect 4632 -1008 4642 -780
rect 4708 -1008 4718 -780
rect 3326 -1072 3388 -1054
rect 3616 -1072 4760 -1068
rect 1856 -1082 3000 -1076
rect 1446 -1134 3000 -1082
rect 1856 -1136 3000 -1134
rect 3326 -1128 4760 -1072
rect 2200 -1238 2210 -1168
rect 2362 -1238 2372 -1168
rect 1318 -1342 1518 -1252
rect 3326 -1304 3388 -1128
rect 3980 -1174 4124 -1172
rect 3980 -1178 4020 -1174
rect 4076 -1178 4124 -1174
rect 3980 -1224 3992 -1178
rect 4112 -1224 4124 -1178
rect 3980 -1226 4020 -1224
rect 4076 -1226 4124 -1224
rect 3980 -1230 4124 -1226
rect 3286 -1342 3390 -1304
rect 1318 -1438 3390 -1342
rect 6550 -1382 6750 -1316
rect 1318 -1452 1518 -1438
rect 6550 -1464 6602 -1382
rect 6700 -1464 6750 -1382
rect 6550 -1516 6750 -1464
rect 2252 -1572 2354 -1566
rect 2252 -1576 2264 -1572
rect 2342 -1576 2354 -1572
rect 3962 -1576 4190 -1572
rect 2218 -1646 2228 -1576
rect 2380 -1646 2390 -1576
rect 3962 -1578 4030 -1576
rect 4108 -1578 4190 -1576
rect 2252 -1650 2264 -1646
rect 2342 -1650 2354 -1646
rect 2252 -1656 2354 -1650
rect 3962 -1648 3974 -1578
rect 4178 -1648 4190 -1578
rect 3962 -1650 4030 -1648
rect 4108 -1650 4190 -1648
rect 3962 -1654 4190 -1650
rect 1848 -1694 4066 -1692
rect 1328 -1750 4756 -1694
rect 1474 -2144 1550 -1750
rect 1848 -1752 4756 -1750
rect 3612 -1754 4756 -1752
rect 1800 -2050 1810 -1838
rect 1868 -2050 1878 -1838
rect 2036 -2038 2046 -1826
rect 2104 -2038 2114 -1826
rect 2270 -2040 2280 -1828
rect 2338 -2040 2348 -1828
rect 2510 -2034 2520 -1822
rect 2578 -2034 2588 -1822
rect 2744 -2032 2754 -1820
rect 2812 -2032 2822 -1820
rect 2980 -2026 2990 -1814
rect 3048 -2026 3058 -1814
rect 3550 -2014 3560 -1824
rect 3636 -2014 3646 -1824
rect 3784 -2004 3794 -1814
rect 3870 -2004 3880 -1814
rect 4020 -1998 4030 -1808
rect 4106 -1998 4116 -1808
rect 4264 -1992 4274 -1802
rect 4350 -1992 4360 -1802
rect 4498 -1994 4508 -1804
rect 4584 -1994 4594 -1804
rect 4730 -1998 4740 -1808
rect 4816 -1998 4826 -1808
rect 1338 -2162 1550 -2144
rect 1338 -2362 1546 -2162
rect 1338 -2366 1550 -2362
rect 1474 -2812 1550 -2366
rect 1914 -2754 1924 -2574
rect 1982 -2754 1992 -2574
rect 2152 -2746 2162 -2566
rect 2220 -2746 2230 -2566
rect 2384 -2754 2394 -2574
rect 2452 -2754 2462 -2574
rect 2622 -2752 2632 -2572
rect 2690 -2752 2700 -2572
rect 2860 -2744 2870 -2564
rect 2928 -2744 2938 -2564
rect 3076 -2596 3538 -2590
rect 3076 -2760 3088 -2596
rect 3526 -2760 3538 -2596
rect 3668 -2760 3678 -2570
rect 3754 -2760 3764 -2570
rect 3904 -2760 3914 -2570
rect 3990 -2760 4000 -2570
rect 4144 -2758 4154 -2568
rect 4230 -2758 4240 -2568
rect 3076 -2766 3538 -2760
rect 4380 -2764 4390 -2574
rect 4466 -2764 4476 -2574
rect 4608 -2766 4618 -2576
rect 4694 -2766 4704 -2576
rect 1472 -2814 2256 -2812
rect 1472 -2824 2982 -2814
rect 1472 -2868 4752 -2824
rect 1474 -2872 1550 -2868
rect 1838 -2874 4752 -2868
rect 2912 -2880 4752 -2874
rect 3608 -2884 4752 -2880
rect 3214 -3204 3414 -3132
rect 3214 -3274 3268 -3204
rect 3352 -3274 3414 -3204
rect 3214 -3332 3414 -3274
<< via1 >>
rect 3270 1866 3352 1952
rect 2678 1672 2864 1684
rect 2678 1624 2710 1672
rect 2710 1624 2840 1672
rect 2840 1624 2864 1672
rect 2678 1610 2864 1624
rect 3624 1688 3820 1708
rect 3624 1626 3652 1688
rect 3652 1626 3796 1688
rect 3796 1626 3820 1688
rect 3624 1616 3820 1626
rect 1816 1244 1876 1448
rect 2052 1252 2112 1456
rect 2286 1248 2346 1452
rect 2524 1252 2584 1456
rect 2760 1260 2820 1464
rect 2998 1266 3058 1470
rect 1918 506 1978 710
rect 2154 512 2214 716
rect 2392 512 2452 716
rect 2630 512 2690 716
rect 3568 1222 3630 1444
rect 3804 1216 3866 1438
rect 4042 1220 4104 1442
rect 4276 1224 4338 1446
rect 4510 1224 4572 1446
rect 4752 1234 4814 1456
rect 2864 508 2924 712
rect 3280 526 3338 712
rect 3694 498 3756 720
rect 3932 504 3994 726
rect 4166 508 4228 730
rect 4398 510 4460 732
rect 4642 510 4704 732
rect 5290 582 5520 610
rect 5290 490 5338 582
rect 5338 490 5484 582
rect 5484 490 5520 582
rect 5290 488 5520 490
rect 5100 126 5178 272
rect 1804 -308 1868 -74
rect 2042 -304 2106 -70
rect 2276 -296 2340 -62
rect 2514 -292 2578 -58
rect 2748 -290 2812 -56
rect 2986 -290 3050 -56
rect 1924 -1034 1988 -800
rect 2158 -1034 2222 -800
rect 2398 -1032 2462 -798
rect 2632 -1032 2696 -798
rect 2870 -1028 2934 -794
rect 3578 -362 3630 -108
rect 3808 -362 3864 -114
rect 4044 -356 4100 -108
rect 4284 -348 4340 -100
rect 4520 -336 4576 -88
rect 4754 -330 4810 -82
rect 5364 100 5432 310
rect 5602 100 5670 310
rect 5846 104 5914 314
rect 6076 104 6144 314
rect 6314 108 6382 318
rect 6546 106 6614 316
rect 5484 -622 5552 -412
rect 5718 -618 5786 -408
rect 5956 -620 6024 -410
rect 6188 -624 6256 -414
rect 6428 -618 6496 -408
rect 3694 -1002 3760 -774
rect 3932 -1000 3998 -772
rect 4170 -1002 4236 -774
rect 4408 -1002 4474 -774
rect 4642 -1008 4708 -780
rect 2210 -1176 2362 -1168
rect 2210 -1228 2234 -1176
rect 2234 -1228 2332 -1176
rect 2332 -1228 2362 -1176
rect 2210 -1238 2362 -1228
rect 4020 -1178 4076 -1174
rect 4020 -1224 4076 -1178
rect 4020 -1226 4076 -1224
rect 6602 -1464 6700 -1382
rect 2228 -1646 2264 -1576
rect 2264 -1646 2342 -1576
rect 2342 -1646 2380 -1576
rect 4030 -1578 4108 -1576
rect 4030 -1648 4108 -1578
rect 4030 -1650 4108 -1648
rect 1810 -2050 1868 -1838
rect 2046 -2038 2104 -1826
rect 2280 -2040 2338 -1828
rect 2520 -2034 2578 -1822
rect 2754 -2032 2812 -1820
rect 2990 -2026 3048 -1814
rect 3560 -2014 3636 -1824
rect 3794 -2004 3870 -1814
rect 4030 -1998 4106 -1808
rect 4274 -1992 4350 -1802
rect 4508 -1994 4584 -1804
rect 4740 -1998 4816 -1808
rect 1924 -2754 1982 -2574
rect 2162 -2746 2220 -2566
rect 2394 -2754 2452 -2574
rect 2632 -2752 2690 -2572
rect 2870 -2744 2928 -2564
rect 3224 -2758 3380 -2626
rect 3678 -2760 3754 -2570
rect 3914 -2760 3990 -2570
rect 4154 -2758 4230 -2568
rect 4390 -2764 4466 -2574
rect 4618 -2766 4694 -2576
rect 3268 -3274 3352 -3204
<< metal2 >>
rect 3270 1952 3352 1962
rect 2724 1866 3270 1950
rect 3352 1866 3796 1950
rect 2724 1854 3796 1866
rect 2728 1694 2818 1854
rect 3684 1718 3770 1854
rect 3624 1708 3820 1718
rect 2678 1684 2864 1694
rect 2678 1600 2864 1610
rect 3624 1606 3820 1616
rect 2728 1474 2818 1600
rect 1816 1448 1876 1458
rect 1798 1266 1816 1446
rect 2052 1456 2112 1466
rect 1876 1266 2052 1446
rect 1816 1234 1876 1244
rect 2286 1452 2346 1462
rect 2112 1266 2286 1446
rect 2052 1242 2112 1252
rect 2524 1456 2584 1466
rect 2346 1266 2524 1446
rect 2286 1238 2346 1248
rect 2728 1464 2820 1474
rect 2728 1446 2760 1464
rect 2584 1266 2760 1446
rect 2524 1242 2584 1252
rect 2998 1470 3058 1480
rect 2820 1266 2998 1446
rect 3568 1452 3630 1454
rect 3684 1452 3770 1606
rect 4752 1456 4814 1466
rect 4276 1452 4338 1456
rect 4510 1452 4572 1456
rect 3556 1446 4752 1452
rect 3058 1266 3076 1446
rect 3556 1444 4276 1446
rect 2760 1250 2820 1260
rect 2998 1256 3058 1266
rect 3556 1232 3568 1444
rect 3630 1442 4276 1444
rect 3630 1438 4042 1442
rect 3630 1232 3804 1438
rect 3568 1212 3630 1222
rect 3866 1232 4042 1438
rect 3804 1206 3866 1216
rect 4104 1232 4276 1442
rect 4042 1210 4104 1220
rect 4338 1232 4510 1446
rect 4276 1214 4338 1224
rect 4572 1234 4752 1446
rect 4814 1234 4828 1452
rect 4572 1232 4828 1234
rect 4752 1224 4814 1232
rect 4510 1214 4572 1224
rect 1918 712 1978 720
rect 2154 716 2214 726
rect 1908 710 2154 712
rect 1908 508 1918 710
rect 1912 506 1918 508
rect 1978 512 2154 710
rect 2392 716 2452 726
rect 2214 512 2392 712
rect 2630 716 2690 726
rect 3694 724 3756 730
rect 3932 726 3994 736
rect 3694 722 3762 724
rect 2452 512 2630 712
rect 2864 712 2924 722
rect 3280 712 3338 722
rect 3678 720 3932 722
rect 2690 512 2864 712
rect 1978 508 2864 512
rect 2924 526 3280 712
rect 3338 526 3346 712
rect 2924 510 3346 526
rect 3678 510 3694 720
rect 2924 508 2940 510
rect 1978 506 1992 508
rect 1804 -74 1868 -64
rect 1782 -286 1804 -76
rect 1912 -76 1992 506
rect 2154 502 2214 508
rect 2392 502 2452 508
rect 2630 502 2690 508
rect 2864 498 2924 508
rect 3756 510 3932 720
rect 3756 498 3762 510
rect 3694 488 3762 498
rect 4166 730 4228 740
rect 3994 510 4166 722
rect 3932 494 3994 504
rect 4398 732 4460 742
rect 4228 510 4398 722
rect 4642 732 4704 742
rect 4460 510 4642 722
rect 4704 510 4718 722
rect 4166 498 4228 508
rect 4398 500 4460 510
rect 2042 -70 2106 -60
rect 1868 -286 2042 -76
rect 1804 -318 1868 -308
rect 2276 -62 2340 -52
rect 2106 -286 2276 -76
rect 2042 -314 2106 -304
rect 2514 -58 2578 -48
rect 2340 -286 2514 -76
rect 2276 -306 2340 -296
rect 2748 -56 2812 -46
rect 2578 -286 2748 -76
rect 2514 -302 2578 -292
rect 2986 -56 3050 -46
rect 2812 -286 2986 -76
rect 2748 -300 2812 -290
rect 3050 -286 3072 -76
rect 3696 -84 3762 488
rect 4620 270 4718 510
rect 5290 610 5520 620
rect 5290 478 5520 488
rect 5398 320 5476 478
rect 5364 312 5476 320
rect 5602 312 5670 320
rect 5846 314 5914 324
rect 5348 310 5846 312
rect 5100 272 5178 282
rect 4618 126 5100 270
rect 4520 -84 4576 -78
rect 4620 -84 4718 126
rect 5100 116 5178 126
rect 5348 104 5364 310
rect 5432 104 5602 310
rect 5364 90 5432 100
rect 5670 104 5846 310
rect 6076 314 6144 324
rect 5914 104 6076 312
rect 6314 318 6382 328
rect 6144 108 6314 312
rect 6546 316 6614 326
rect 6382 108 6546 312
rect 6144 106 6546 108
rect 6614 106 6628 312
rect 6144 104 6628 106
rect 5602 90 5670 100
rect 5846 94 5914 104
rect 6076 94 6144 104
rect 6314 98 6382 104
rect 6546 96 6614 104
rect 4754 -82 4810 -72
rect 3560 -88 4754 -84
rect 3560 -100 4520 -88
rect 3560 -108 4284 -100
rect 2986 -300 3050 -290
rect 3560 -362 3578 -108
rect 3630 -114 4044 -108
rect 3630 -362 3808 -114
rect 3864 -356 4044 -114
rect 4100 -348 4284 -108
rect 4340 -336 4520 -100
rect 4576 -330 4754 -88
rect 4810 -330 4830 -84
rect 4576 -336 4830 -330
rect 4340 -348 4830 -336
rect 4100 -356 4830 -348
rect 3864 -362 4830 -356
rect 3560 -364 4830 -362
rect 3578 -372 3630 -364
rect 3808 -372 3864 -364
rect 4044 -366 4100 -364
rect 5484 -412 5552 -402
rect 5464 -618 5484 -420
rect 5718 -408 5786 -398
rect 5552 -618 5718 -420
rect 5956 -410 6024 -400
rect 5786 -618 5956 -420
rect 5484 -632 5552 -622
rect 3694 -774 3760 -764
rect 1924 -798 1988 -790
rect 2158 -798 2222 -790
rect 2398 -798 2462 -788
rect 2632 -798 2696 -788
rect 2870 -794 2934 -784
rect 1902 -800 2398 -798
rect 1902 -1026 1924 -800
rect 1920 -1034 1924 -1026
rect 1988 -1026 2158 -800
rect 1988 -1034 1994 -1026
rect 1810 -1838 1868 -1828
rect 1780 -2024 1810 -1840
rect 1920 -1840 1994 -1034
rect 2222 -1026 2398 -800
rect 2158 -1044 2222 -1034
rect 2462 -1026 2632 -798
rect 2398 -1042 2462 -1032
rect 2696 -1026 2870 -798
rect 2632 -1042 2696 -1032
rect 2934 -858 2956 -798
rect 3676 -858 3694 -776
rect 2934 -946 3694 -858
rect 2934 -1026 2956 -946
rect 3676 -1002 3694 -946
rect 3932 -772 3998 -762
rect 3760 -1000 3932 -776
rect 4170 -774 4236 -764
rect 3998 -1000 4170 -776
rect 3760 -1002 4170 -1000
rect 4408 -774 4474 -764
rect 4236 -1002 4408 -776
rect 4642 -776 4708 -770
rect 4474 -780 4722 -776
rect 4474 -1002 4642 -780
rect 3676 -1008 4642 -1002
rect 4708 -1008 4722 -780
rect 3676 -1012 4722 -1008
rect 4642 -1018 4708 -1012
rect 2870 -1038 2934 -1028
rect 2210 -1168 2362 -1158
rect 4020 -1172 4076 -1164
rect 2210 -1248 2362 -1238
rect 4008 -1174 4104 -1172
rect 4008 -1226 4020 -1174
rect 4076 -1226 4104 -1174
rect 5596 -1182 5670 -618
rect 5718 -628 5786 -618
rect 6188 -414 6256 -404
rect 6024 -618 6188 -420
rect 5956 -630 6024 -620
rect 6428 -408 6496 -398
rect 6256 -618 6428 -420
rect 6496 -618 6510 -420
rect 6188 -634 6256 -624
rect 6428 -628 6496 -618
rect 2254 -1566 2336 -1248
rect 4008 -1566 4104 -1226
rect 5594 -1198 5670 -1182
rect 5594 -1360 5668 -1198
rect 5594 -1382 6700 -1360
rect 5594 -1464 6602 -1382
rect 5594 -1482 6700 -1464
rect 2228 -1576 2380 -1566
rect 2228 -1656 2380 -1646
rect 4008 -1576 4108 -1566
rect 4008 -1650 4030 -1576
rect 4008 -1654 4108 -1650
rect 4030 -1660 4108 -1654
rect 5594 -1790 5668 -1482
rect 2046 -1826 2104 -1816
rect 1868 -2024 2046 -1840
rect 2280 -1828 2338 -1818
rect 2104 -2024 2280 -1840
rect 2046 -2048 2104 -2038
rect 2520 -1822 2578 -1812
rect 2338 -2024 2520 -1840
rect 2280 -2050 2338 -2040
rect 2754 -1820 2812 -1810
rect 2578 -2024 2754 -1840
rect 2520 -2044 2578 -2034
rect 2990 -1814 3048 -1804
rect 3794 -1814 3870 -1804
rect 2812 -2024 2990 -1840
rect 2754 -2042 2812 -2032
rect 3560 -1816 3636 -1814
rect 3536 -1824 3794 -1816
rect 3048 -2024 3068 -1840
rect 3536 -2002 3560 -1824
rect 3636 -2002 3794 -1824
rect 4030 -1808 4106 -1798
rect 3870 -1998 4030 -1816
rect 4274 -1802 4350 -1792
rect 4106 -1992 4274 -1816
rect 4508 -1804 4584 -1794
rect 4350 -1992 4508 -1816
rect 4106 -1994 4508 -1992
rect 4740 -1808 4816 -1798
rect 4584 -1994 4740 -1816
rect 4106 -1998 4740 -1994
rect 4816 -1856 4822 -1816
rect 5596 -1854 5666 -1790
rect 5064 -1856 5672 -1854
rect 4816 -1928 5672 -1856
rect 4816 -1930 5348 -1928
rect 4816 -1998 4822 -1930
rect 5596 -1934 5666 -1928
rect 3870 -2002 4822 -1998
rect 3794 -2014 3870 -2004
rect 4030 -2008 4106 -2002
rect 4508 -2004 4584 -2002
rect 4740 -2008 4816 -2002
rect 3560 -2024 3636 -2014
rect 2990 -2036 3048 -2026
rect 1810 -2060 1868 -2050
rect 1924 -2574 1982 -2564
rect 1906 -2746 1924 -2578
rect 2162 -2566 2220 -2556
rect 1982 -2746 2162 -2578
rect 2394 -2574 2452 -2564
rect 2220 -2746 2394 -2578
rect 1924 -2764 1982 -2754
rect 2162 -2756 2220 -2746
rect 2632 -2572 2690 -2562
rect 2452 -2746 2632 -2578
rect 2394 -2764 2452 -2754
rect 2870 -2564 2928 -2554
rect 2690 -2744 2870 -2578
rect 3678 -2570 3754 -2560
rect 2928 -2640 2940 -2578
rect 3228 -2616 3386 -2614
rect 3224 -2626 3386 -2616
rect 2928 -2724 3224 -2640
rect 2928 -2744 2940 -2724
rect 2690 -2746 2940 -2744
rect 2632 -2762 2690 -2752
rect 2870 -2754 2928 -2746
rect 3380 -2640 3386 -2626
rect 3664 -2640 3678 -2574
rect 3380 -2724 3678 -2640
rect 3380 -2758 3386 -2724
rect 3224 -2768 3386 -2758
rect 3664 -2760 3678 -2724
rect 3914 -2570 3990 -2560
rect 3754 -2760 3914 -2574
rect 4154 -2568 4230 -2558
rect 3990 -2758 4154 -2574
rect 4390 -2574 4466 -2564
rect 4618 -2574 4694 -2566
rect 4230 -2758 4390 -2574
rect 3990 -2760 4390 -2758
rect 3664 -2762 4390 -2760
rect 3228 -3204 3386 -2768
rect 3678 -2770 3754 -2762
rect 3914 -2770 3990 -2762
rect 4154 -2768 4230 -2762
rect 4466 -2576 4694 -2574
rect 4466 -2762 4618 -2576
rect 4390 -2774 4466 -2764
rect 4618 -2776 4694 -2766
rect 3228 -3274 3268 -3204
rect 3352 -3274 3386 -3204
rect 3228 -3282 3386 -3274
rect 3268 -3284 3352 -3282
use sky130_fd_pr__nfet_01v8_4H4H2H  XM1
timestamp 1706794580
transform 1 0 2427 0 1 -546
box -757 -710 757 710
use sky130_fd_pr__nfet_01v8_4H4H2H  XM2
timestamp 1706794580
transform 1 0 4197 0 1 -540
box -757 -710 757 710
use sky130_fd_pr__pfet_01v8_4C76A3  XM3
timestamp 1706798884
transform 1 0 2423 0 1 977
box -757 -719 757 719
use sky130_fd_pr__pfet_01v8_4C76A3  XM4
timestamp 1706798884
transform 1 0 4197 0 1 981
box -757 -719 757 719
use sky130_fd_pr__nfet_01v8_4H4H2H  XM5
timestamp 1706794580
transform 1 0 2425 0 1 -2284
box -757 -710 757 710
use sky130_fd_pr__pfet_01v8_4C76A3  XM6
timestamp 1706798884
transform 1 0 5987 0 1 -145
box -757 -719 757 719
use sky130_fd_pr__nfet_01v8_4H4H2H  XM7
timestamp 1706794580
transform 1 0 4189 0 1 -2290
box -757 -710 757 710
<< labels >>
flabel metal1 1288 -668 1488 -468 0 FreeSans 256 0 0 0 inp1
port 0 nsew
flabel metal1 1318 -1452 1518 -1252 0 FreeSans 256 0 0 0 inp2
port 1 nsew
flabel metal1 1338 -2366 1546 -2144 0 FreeSans 1600 0 0 0 vbias
port 7 nsew
flabel metal1 6550 -1516 6750 -1316 0 FreeSans 256 0 0 0 vout
port 5 nsew
flabel metal1 3210 1808 3410 2008 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 3214 -3332 3414 -3132 0 FreeSans 256 0 0 0 vss
port 3 nsew
<< end >>
