magic
tech sky130A
magscale 1 2
timestamp 1706788245
<< error_p >>
rect -560 572 -502 578
rect -442 572 -384 578
rect -324 572 -266 578
rect -206 572 -148 578
rect -88 572 -30 578
rect 30 572 88 578
rect 148 572 206 578
rect 266 572 324 578
rect 384 572 442 578
rect 502 572 560 578
rect -560 538 -548 572
rect -442 538 -430 572
rect -324 538 -312 572
rect -206 538 -194 572
rect -88 538 -76 572
rect 30 538 42 572
rect 148 538 160 572
rect 266 538 278 572
rect 384 538 396 572
rect 502 538 514 572
rect -560 532 -502 538
rect -442 532 -384 538
rect -324 532 -266 538
rect -206 532 -148 538
rect -88 532 -30 538
rect 30 532 88 538
rect 148 532 206 538
rect 266 532 324 538
rect 384 532 442 538
rect 502 532 560 538
rect -560 -538 -502 -532
rect -442 -538 -384 -532
rect -324 -538 -266 -532
rect -206 -538 -148 -532
rect -88 -538 -30 -532
rect 30 -538 88 -532
rect 148 -538 206 -532
rect 266 -538 324 -532
rect 384 -538 442 -532
rect 502 -538 560 -532
rect -560 -572 -548 -538
rect -442 -572 -430 -538
rect -324 -572 -312 -538
rect -206 -572 -194 -538
rect -88 -572 -76 -538
rect 30 -572 42 -538
rect 148 -572 160 -538
rect 266 -572 278 -538
rect 384 -572 396 -538
rect 502 -572 514 -538
rect -560 -578 -502 -572
rect -442 -578 -384 -572
rect -324 -578 -266 -572
rect -206 -578 -148 -572
rect -88 -578 -30 -572
rect 30 -578 88 -572
rect 148 -578 206 -572
rect 266 -578 324 -572
rect 384 -578 442 -572
rect 502 -578 560 -572
<< pwell >>
rect -757 -710 757 710
<< nmos >>
rect -561 -500 -501 500
rect -443 -500 -383 500
rect -325 -500 -265 500
rect -207 -500 -147 500
rect -89 -500 -29 500
rect 29 -500 89 500
rect 147 -500 207 500
rect 265 -500 325 500
rect 383 -500 443 500
rect 501 -500 561 500
<< ndiff >>
rect -619 488 -561 500
rect -619 -488 -607 488
rect -573 -488 -561 488
rect -619 -500 -561 -488
rect -501 488 -443 500
rect -501 -488 -489 488
rect -455 -488 -443 488
rect -501 -500 -443 -488
rect -383 488 -325 500
rect -383 -488 -371 488
rect -337 -488 -325 488
rect -383 -500 -325 -488
rect -265 488 -207 500
rect -265 -488 -253 488
rect -219 -488 -207 488
rect -265 -500 -207 -488
rect -147 488 -89 500
rect -147 -488 -135 488
rect -101 -488 -89 488
rect -147 -500 -89 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 89 488 147 500
rect 89 -488 101 488
rect 135 -488 147 488
rect 89 -500 147 -488
rect 207 488 265 500
rect 207 -488 219 488
rect 253 -488 265 488
rect 207 -500 265 -488
rect 325 488 383 500
rect 325 -488 337 488
rect 371 -488 383 488
rect 325 -500 383 -488
rect 443 488 501 500
rect 443 -488 455 488
rect 489 -488 501 488
rect 443 -500 501 -488
rect 561 488 619 500
rect 561 -488 573 488
rect 607 -488 619 488
rect 561 -500 619 -488
<< ndiffc >>
rect -607 -488 -573 488
rect -489 -488 -455 488
rect -371 -488 -337 488
rect -253 -488 -219 488
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
rect 219 -488 253 488
rect 337 -488 371 488
rect 455 -488 489 488
rect 573 -488 607 488
<< psubdiff >>
rect -721 640 -625 674
rect 625 640 721 674
rect -721 578 -687 640
rect 687 578 721 640
rect -721 -640 -687 -578
rect 687 -640 721 -578
rect -721 -674 -625 -640
rect 625 -674 721 -640
<< psubdiffcont >>
rect -625 640 625 674
rect -721 -578 -687 578
rect 687 -578 721 578
rect -625 -674 625 -640
<< poly >>
rect -564 572 -498 588
rect -564 538 -548 572
rect -514 538 -498 572
rect -564 522 -498 538
rect -446 572 -380 588
rect -446 538 -430 572
rect -396 538 -380 572
rect -446 522 -380 538
rect -328 572 -262 588
rect -328 538 -312 572
rect -278 538 -262 572
rect -328 522 -262 538
rect -210 572 -144 588
rect -210 538 -194 572
rect -160 538 -144 572
rect -210 522 -144 538
rect -92 572 -26 588
rect -92 538 -76 572
rect -42 538 -26 572
rect -92 522 -26 538
rect 26 572 92 588
rect 26 538 42 572
rect 76 538 92 572
rect 26 522 92 538
rect 144 572 210 588
rect 144 538 160 572
rect 194 538 210 572
rect 144 522 210 538
rect 262 572 328 588
rect 262 538 278 572
rect 312 538 328 572
rect 262 522 328 538
rect 380 572 446 588
rect 380 538 396 572
rect 430 538 446 572
rect 380 522 446 538
rect 498 572 564 588
rect 498 538 514 572
rect 548 538 564 572
rect 498 522 564 538
rect -561 500 -501 522
rect -443 500 -383 522
rect -325 500 -265 522
rect -207 500 -147 522
rect -89 500 -29 522
rect 29 500 89 522
rect 147 500 207 522
rect 265 500 325 522
rect 383 500 443 522
rect 501 500 561 522
rect -561 -522 -501 -500
rect -443 -522 -383 -500
rect -325 -522 -265 -500
rect -207 -522 -147 -500
rect -89 -522 -29 -500
rect 29 -522 89 -500
rect 147 -522 207 -500
rect 265 -522 325 -500
rect 383 -522 443 -500
rect 501 -522 561 -500
rect -564 -538 -498 -522
rect -564 -572 -548 -538
rect -514 -572 -498 -538
rect -564 -588 -498 -572
rect -446 -538 -380 -522
rect -446 -572 -430 -538
rect -396 -572 -380 -538
rect -446 -588 -380 -572
rect -328 -538 -262 -522
rect -328 -572 -312 -538
rect -278 -572 -262 -538
rect -328 -588 -262 -572
rect -210 -538 -144 -522
rect -210 -572 -194 -538
rect -160 -572 -144 -538
rect -210 -588 -144 -572
rect -92 -538 -26 -522
rect -92 -572 -76 -538
rect -42 -572 -26 -538
rect -92 -588 -26 -572
rect 26 -538 92 -522
rect 26 -572 42 -538
rect 76 -572 92 -538
rect 26 -588 92 -572
rect 144 -538 210 -522
rect 144 -572 160 -538
rect 194 -572 210 -538
rect 144 -588 210 -572
rect 262 -538 328 -522
rect 262 -572 278 -538
rect 312 -572 328 -538
rect 262 -588 328 -572
rect 380 -538 446 -522
rect 380 -572 396 -538
rect 430 -572 446 -538
rect 380 -588 446 -572
rect 498 -538 564 -522
rect 498 -572 514 -538
rect 548 -572 564 -538
rect 498 -588 564 -572
<< polycont >>
rect -548 538 -514 572
rect -430 538 -396 572
rect -312 538 -278 572
rect -194 538 -160 572
rect -76 538 -42 572
rect 42 538 76 572
rect 160 538 194 572
rect 278 538 312 572
rect 396 538 430 572
rect 514 538 548 572
rect -548 -572 -514 -538
rect -430 -572 -396 -538
rect -312 -572 -278 -538
rect -194 -572 -160 -538
rect -76 -572 -42 -538
rect 42 -572 76 -538
rect 160 -572 194 -538
rect 278 -572 312 -538
rect 396 -572 430 -538
rect 514 -572 548 -538
<< locali >>
rect -721 640 -625 674
rect 625 640 721 674
rect -721 578 -687 640
rect 687 578 721 640
rect -564 538 -548 572
rect -514 538 -498 572
rect -446 538 -430 572
rect -396 538 -380 572
rect -328 538 -312 572
rect -278 538 -262 572
rect -210 538 -194 572
rect -160 538 -144 572
rect -92 538 -76 572
rect -42 538 -26 572
rect 26 538 42 572
rect 76 538 92 572
rect 144 538 160 572
rect 194 538 210 572
rect 262 538 278 572
rect 312 538 328 572
rect 380 538 396 572
rect 430 538 446 572
rect 498 538 514 572
rect 548 538 564 572
rect -607 488 -573 504
rect -607 -504 -573 -488
rect -489 488 -455 504
rect -489 -504 -455 -488
rect -371 488 -337 504
rect -371 -504 -337 -488
rect -253 488 -219 504
rect -253 -504 -219 -488
rect -135 488 -101 504
rect -135 -504 -101 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 101 488 135 504
rect 101 -504 135 -488
rect 219 488 253 504
rect 219 -504 253 -488
rect 337 488 371 504
rect 337 -504 371 -488
rect 455 488 489 504
rect 455 -504 489 -488
rect 573 488 607 504
rect 573 -504 607 -488
rect -564 -572 -548 -538
rect -514 -572 -498 -538
rect -446 -572 -430 -538
rect -396 -572 -380 -538
rect -328 -572 -312 -538
rect -278 -572 -262 -538
rect -210 -572 -194 -538
rect -160 -572 -144 -538
rect -92 -572 -76 -538
rect -42 -572 -26 -538
rect 26 -572 42 -538
rect 76 -572 92 -538
rect 144 -572 160 -538
rect 194 -572 210 -538
rect 262 -572 278 -538
rect 312 -572 328 -538
rect 380 -572 396 -538
rect 430 -572 446 -538
rect 498 -572 514 -538
rect 548 -572 564 -538
rect -721 -640 -687 -578
rect 687 -640 721 -578
rect -721 -674 -625 -640
rect 625 -674 721 -640
<< viali >>
rect -548 538 -514 572
rect -430 538 -396 572
rect -312 538 -278 572
rect -194 538 -160 572
rect -76 538 -42 572
rect 42 538 76 572
rect 160 538 194 572
rect 278 538 312 572
rect 396 538 430 572
rect 514 538 548 572
rect -607 -488 -573 488
rect -489 -488 -455 488
rect -371 -488 -337 488
rect -253 -488 -219 488
rect -135 -488 -101 488
rect -17 -488 17 488
rect 101 -488 135 488
rect 219 -488 253 488
rect 337 -488 371 488
rect 455 -488 489 488
rect 573 -488 607 488
rect -548 -572 -514 -538
rect -430 -572 -396 -538
rect -312 -572 -278 -538
rect -194 -572 -160 -538
rect -76 -572 -42 -538
rect 42 -572 76 -538
rect 160 -572 194 -538
rect 278 -572 312 -538
rect 396 -572 430 -538
rect 514 -572 548 -538
<< metal1 >>
rect -560 572 -502 578
rect -560 538 -548 572
rect -514 538 -502 572
rect -560 532 -502 538
rect -442 572 -384 578
rect -442 538 -430 572
rect -396 538 -384 572
rect -442 532 -384 538
rect -324 572 -266 578
rect -324 538 -312 572
rect -278 538 -266 572
rect -324 532 -266 538
rect -206 572 -148 578
rect -206 538 -194 572
rect -160 538 -148 572
rect -206 532 -148 538
rect -88 572 -30 578
rect -88 538 -76 572
rect -42 538 -30 572
rect -88 532 -30 538
rect 30 572 88 578
rect 30 538 42 572
rect 76 538 88 572
rect 30 532 88 538
rect 148 572 206 578
rect 148 538 160 572
rect 194 538 206 572
rect 148 532 206 538
rect 266 572 324 578
rect 266 538 278 572
rect 312 538 324 572
rect 266 532 324 538
rect 384 572 442 578
rect 384 538 396 572
rect 430 538 442 572
rect 384 532 442 538
rect 502 572 560 578
rect 502 538 514 572
rect 548 538 560 572
rect 502 532 560 538
rect -613 488 -567 500
rect -613 -488 -607 488
rect -573 -488 -567 488
rect -613 -500 -567 -488
rect -495 488 -449 500
rect -495 -488 -489 488
rect -455 -488 -449 488
rect -495 -500 -449 -488
rect -377 488 -331 500
rect -377 -488 -371 488
rect -337 -488 -331 488
rect -377 -500 -331 -488
rect -259 488 -213 500
rect -259 -488 -253 488
rect -219 -488 -213 488
rect -259 -500 -213 -488
rect -141 488 -95 500
rect -141 -488 -135 488
rect -101 -488 -95 488
rect -141 -500 -95 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 95 488 141 500
rect 95 -488 101 488
rect 135 -488 141 488
rect 95 -500 141 -488
rect 213 488 259 500
rect 213 -488 219 488
rect 253 -488 259 488
rect 213 -500 259 -488
rect 331 488 377 500
rect 331 -488 337 488
rect 371 -488 377 488
rect 331 -500 377 -488
rect 449 488 495 500
rect 449 -488 455 488
rect 489 -488 495 488
rect 449 -500 495 -488
rect 567 488 613 500
rect 567 -488 573 488
rect 607 -488 613 488
rect 567 -500 613 -488
rect -560 -538 -502 -532
rect -560 -572 -548 -538
rect -514 -572 -502 -538
rect -560 -578 -502 -572
rect -442 -538 -384 -532
rect -442 -572 -430 -538
rect -396 -572 -384 -538
rect -442 -578 -384 -572
rect -324 -538 -266 -532
rect -324 -572 -312 -538
rect -278 -572 -266 -538
rect -324 -578 -266 -572
rect -206 -538 -148 -532
rect -206 -572 -194 -538
rect -160 -572 -148 -538
rect -206 -578 -148 -572
rect -88 -538 -30 -532
rect -88 -572 -76 -538
rect -42 -572 -30 -538
rect -88 -578 -30 -572
rect 30 -538 88 -532
rect 30 -572 42 -538
rect 76 -572 88 -538
rect 30 -578 88 -572
rect 148 -538 206 -532
rect 148 -572 160 -538
rect 194 -572 206 -538
rect 148 -578 206 -572
rect 266 -538 324 -532
rect 266 -572 278 -538
rect 312 -572 324 -538
rect 266 -578 324 -572
rect 384 -538 442 -532
rect 384 -572 396 -538
rect 430 -572 442 -538
rect 384 -578 442 -572
rect 502 -538 560 -532
rect 502 -572 514 -538
rect 548 -572 560 -538
rect 502 -578 560 -572
<< properties >>
string FIXED_BBOX -704 -657 704 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.300 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
