magic
tech sky130A
magscale 1 2
timestamp 1708951863
<< locali >>
rect -1442 1172 -1432 1216
rect -1430 780 -1396 978
rect -1430 742 -1364 780
rect -1430 736 -80 742
rect -1430 706 -48 736
<< viali >>
rect -1804 1178 -1754 1220
rect -1432 1172 -1398 1216
<< metal1 >>
rect -2468 2178 -1232 2180
rect -2468 2116 -1204 2178
rect -1266 1990 -1204 2116
rect -1430 1832 -1258 1876
rect -1992 1220 -1946 1710
rect -1430 1492 -1398 1832
rect -1816 1220 -1742 1226
rect -1992 1178 -1804 1220
rect -1754 1178 -1742 1220
rect -1992 1176 -1742 1178
rect -1992 1172 -1946 1176
rect -1816 1172 -1742 1176
rect -1444 1218 -1376 1222
rect -1236 1218 -1186 1220
rect -1444 1216 -1186 1218
rect -1444 1172 -1432 1216
rect -1398 1174 -1186 1216
rect -1398 1172 -1376 1174
rect -1444 1166 -1376 1172
rect -1236 1014 -1186 1174
rect -2104 914 -1800 960
rect -1876 446 -1260 484
rect -1876 372 -1828 446
use cp_schem  cp_schem_0
timestamp 1708951863
transform 1 0 -2570 0 1 -3580
box 1298 4024 6324 5767
use pfd  pfd_0
timestamp 1708936645
transform 1 0 -5782 0 1 1874
box 786 -1880 3956 334
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform 1 0 -1826 0 1 962
box -38 -48 498 592
<< end >>
