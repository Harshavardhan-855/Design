** sch_path: /home/harsh/design/xschem/cs_amplifier_tb.sch
.subckt cs_amplifier_tb

x1 net1 output input GND cs_amplifier
V1 input GND sin(0.9 10m 1e6 0)
V2 net1 GND 1.8
C1 output GND 2p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.control
 save all
 tran 0.01u 10u
 write cs_amplifier_tb.raw
 plot v(input) v(output)
.endc


**** end user architecture code
.ends

* expanding   symbol:  cs_amplifier.sym # of pins=4
** sym_path: /home/harsh/design/xschem/cs_amplifier.sym
** sch_path: /home/harsh/design/xschem/cs_amplifier.sch
.subckt cs_amplifier vdd output input gnd
*.PININFO input:I vdd:B gnd:B output:O
XM1 output input gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XR1 output vdd gnd sky130_fd_pr__res_high_po W=1.012 L=2 mult=1 m=1
.ends

.GLOBAL GND
.end
