magic
tech sky130A
magscale 1 2
timestamp 1708941600
<< error_p >>
rect -365 132 -307 138
rect -173 132 -115 138
rect 19 132 77 138
rect 211 132 269 138
rect 403 132 461 138
rect -365 98 -353 132
rect -173 98 -161 132
rect 19 98 31 132
rect 211 98 223 132
rect 403 98 415 132
rect -365 92 -307 98
rect -173 92 -115 98
rect 19 92 77 98
rect 211 92 269 98
rect 403 92 461 98
rect -461 -98 -403 -92
rect -269 -98 -211 -92
rect -77 -98 -19 -92
rect 115 -98 173 -92
rect 307 -98 365 -92
rect -461 -132 -449 -98
rect -269 -132 -257 -98
rect -77 -132 -65 -98
rect 115 -132 127 -98
rect 307 -132 319 -98
rect -461 -138 -403 -132
rect -269 -138 -211 -132
rect -77 -138 -19 -132
rect 115 -138 173 -132
rect 307 -138 365 -132
<< pwell >>
rect -647 -270 647 270
<< nmos >>
rect -447 -60 -417 60
rect -351 -60 -321 60
rect -255 -60 -225 60
rect -159 -60 -129 60
rect -63 -60 -33 60
rect 33 -60 63 60
rect 129 -60 159 60
rect 225 -60 255 60
rect 321 -60 351 60
rect 417 -60 447 60
<< ndiff >>
rect -509 48 -447 60
rect -509 -48 -497 48
rect -463 -48 -447 48
rect -509 -60 -447 -48
rect -417 48 -351 60
rect -417 -48 -401 48
rect -367 -48 -351 48
rect -417 -60 -351 -48
rect -321 48 -255 60
rect -321 -48 -305 48
rect -271 -48 -255 48
rect -321 -60 -255 -48
rect -225 48 -159 60
rect -225 -48 -209 48
rect -175 -48 -159 48
rect -225 -60 -159 -48
rect -129 48 -63 60
rect -129 -48 -113 48
rect -79 -48 -63 48
rect -129 -60 -63 -48
rect -33 48 33 60
rect -33 -48 -17 48
rect 17 -48 33 48
rect -33 -60 33 -48
rect 63 48 129 60
rect 63 -48 79 48
rect 113 -48 129 48
rect 63 -60 129 -48
rect 159 48 225 60
rect 159 -48 175 48
rect 209 -48 225 48
rect 159 -60 225 -48
rect 255 48 321 60
rect 255 -48 271 48
rect 305 -48 321 48
rect 255 -60 321 -48
rect 351 48 417 60
rect 351 -48 367 48
rect 401 -48 417 48
rect 351 -60 417 -48
rect 447 48 509 60
rect 447 -48 463 48
rect 497 -48 509 48
rect 447 -60 509 -48
<< ndiffc >>
rect -497 -48 -463 48
rect -401 -48 -367 48
rect -305 -48 -271 48
rect -209 -48 -175 48
rect -113 -48 -79 48
rect -17 -48 17 48
rect 79 -48 113 48
rect 175 -48 209 48
rect 271 -48 305 48
rect 367 -48 401 48
rect 463 -48 497 48
<< psubdiff >>
rect -611 200 -515 234
rect 515 200 611 234
rect -611 138 -577 200
rect 577 138 611 200
rect -611 -200 -577 -138
rect 577 -200 611 -138
rect -611 -234 -515 -200
rect 515 -234 611 -200
<< psubdiffcont >>
rect -515 200 515 234
rect -611 -138 -577 138
rect 577 -138 611 138
rect -515 -234 515 -200
<< poly >>
rect -369 132 -303 148
rect -369 98 -353 132
rect -319 98 -303 132
rect -447 60 -417 86
rect -369 82 -303 98
rect -177 132 -111 148
rect -177 98 -161 132
rect -127 98 -111 132
rect -351 60 -321 82
rect -255 60 -225 86
rect -177 82 -111 98
rect 15 132 81 148
rect 15 98 31 132
rect 65 98 81 132
rect -159 60 -129 82
rect -63 60 -33 86
rect 15 82 81 98
rect 207 132 273 148
rect 207 98 223 132
rect 257 98 273 132
rect 33 60 63 82
rect 129 60 159 86
rect 207 82 273 98
rect 399 132 465 148
rect 399 98 415 132
rect 449 98 465 132
rect 225 60 255 82
rect 321 60 351 86
rect 399 82 465 98
rect 417 60 447 82
rect -447 -82 -417 -60
rect -465 -98 -399 -82
rect -351 -86 -321 -60
rect -255 -82 -225 -60
rect -465 -132 -449 -98
rect -415 -132 -399 -98
rect -465 -148 -399 -132
rect -273 -98 -207 -82
rect -159 -86 -129 -60
rect -63 -82 -33 -60
rect -273 -132 -257 -98
rect -223 -132 -207 -98
rect -273 -148 -207 -132
rect -81 -98 -15 -82
rect 33 -86 63 -60
rect 129 -82 159 -60
rect -81 -132 -65 -98
rect -31 -132 -15 -98
rect -81 -148 -15 -132
rect 111 -98 177 -82
rect 225 -86 255 -60
rect 321 -82 351 -60
rect 111 -132 127 -98
rect 161 -132 177 -98
rect 111 -148 177 -132
rect 303 -98 369 -82
rect 417 -86 447 -60
rect 303 -132 319 -98
rect 353 -132 369 -98
rect 303 -148 369 -132
<< polycont >>
rect -353 98 -319 132
rect -161 98 -127 132
rect 31 98 65 132
rect 223 98 257 132
rect 415 98 449 132
rect -449 -132 -415 -98
rect -257 -132 -223 -98
rect -65 -132 -31 -98
rect 127 -132 161 -98
rect 319 -132 353 -98
<< locali >>
rect -611 200 -515 234
rect 515 200 611 234
rect -611 138 -577 200
rect 577 138 611 200
rect -369 98 -353 132
rect -319 98 -303 132
rect -177 98 -161 132
rect -127 98 -111 132
rect 15 98 31 132
rect 65 98 81 132
rect 207 98 223 132
rect 257 98 273 132
rect 399 98 415 132
rect 449 98 465 132
rect -497 48 -463 64
rect -497 -64 -463 -48
rect -401 48 -367 64
rect -401 -64 -367 -48
rect -305 48 -271 64
rect -305 -64 -271 -48
rect -209 48 -175 64
rect -209 -64 -175 -48
rect -113 48 -79 64
rect -113 -64 -79 -48
rect -17 48 17 64
rect -17 -64 17 -48
rect 79 48 113 64
rect 79 -64 113 -48
rect 175 48 209 64
rect 175 -64 209 -48
rect 271 48 305 64
rect 271 -64 305 -48
rect 367 48 401 64
rect 367 -64 401 -48
rect 463 48 497 64
rect 463 -64 497 -48
rect -465 -132 -449 -98
rect -415 -132 -399 -98
rect -273 -132 -257 -98
rect -223 -132 -207 -98
rect -81 -132 -65 -98
rect -31 -132 -15 -98
rect 111 -132 127 -98
rect 161 -132 177 -98
rect 303 -132 319 -98
rect 353 -132 369 -98
rect -611 -200 -577 -138
rect 577 -200 611 -138
rect -611 -234 -515 -200
rect 515 -234 611 -200
<< viali >>
rect -353 98 -319 132
rect -161 98 -127 132
rect 31 98 65 132
rect 223 98 257 132
rect 415 98 449 132
rect -497 -48 -463 48
rect -401 -48 -367 48
rect -305 -48 -271 48
rect -209 -48 -175 48
rect -113 -48 -79 48
rect -17 -48 17 48
rect 79 -48 113 48
rect 175 -48 209 48
rect 271 -48 305 48
rect 367 -48 401 48
rect 463 -48 497 48
rect -449 -132 -415 -98
rect -257 -132 -223 -98
rect -65 -132 -31 -98
rect 127 -132 161 -98
rect 319 -132 353 -98
<< metal1 >>
rect -365 132 -307 138
rect -365 98 -353 132
rect -319 98 -307 132
rect -365 92 -307 98
rect -173 132 -115 138
rect -173 98 -161 132
rect -127 98 -115 132
rect -173 92 -115 98
rect 19 132 77 138
rect 19 98 31 132
rect 65 98 77 132
rect 19 92 77 98
rect 211 132 269 138
rect 211 98 223 132
rect 257 98 269 132
rect 211 92 269 98
rect 403 132 461 138
rect 403 98 415 132
rect 449 98 461 132
rect 403 92 461 98
rect -503 48 -457 60
rect -503 -48 -497 48
rect -463 -48 -457 48
rect -503 -60 -457 -48
rect -407 48 -361 60
rect -407 -48 -401 48
rect -367 -48 -361 48
rect -407 -60 -361 -48
rect -311 48 -265 60
rect -311 -48 -305 48
rect -271 -48 -265 48
rect -311 -60 -265 -48
rect -215 48 -169 60
rect -215 -48 -209 48
rect -175 -48 -169 48
rect -215 -60 -169 -48
rect -119 48 -73 60
rect -119 -48 -113 48
rect -79 -48 -73 48
rect -119 -60 -73 -48
rect -23 48 23 60
rect -23 -48 -17 48
rect 17 -48 23 48
rect -23 -60 23 -48
rect 73 48 119 60
rect 73 -48 79 48
rect 113 -48 119 48
rect 73 -60 119 -48
rect 169 48 215 60
rect 169 -48 175 48
rect 209 -48 215 48
rect 169 -60 215 -48
rect 265 48 311 60
rect 265 -48 271 48
rect 305 -48 311 48
rect 265 -60 311 -48
rect 361 48 407 60
rect 361 -48 367 48
rect 401 -48 407 48
rect 361 -60 407 -48
rect 457 48 503 60
rect 457 -48 463 48
rect 497 -48 503 48
rect 457 -60 503 -48
rect -461 -98 -403 -92
rect -461 -132 -449 -98
rect -415 -132 -403 -98
rect -461 -138 -403 -132
rect -269 -98 -211 -92
rect -269 -132 -257 -98
rect -223 -132 -211 -98
rect -269 -138 -211 -132
rect -77 -98 -19 -92
rect -77 -132 -65 -98
rect -31 -132 -19 -98
rect -77 -138 -19 -132
rect 115 -98 173 -92
rect 115 -132 127 -98
rect 161 -132 173 -98
rect 115 -138 173 -132
rect 307 -98 365 -92
rect 307 -132 319 -98
rect 353 -132 365 -98
rect 307 -138 365 -132
<< properties >>
string FIXED_BBOX -594 -217 594 217
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.6 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
