magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -845 372 -787 378
rect -653 372 -595 378
rect -461 372 -403 378
rect -269 372 -211 378
rect -77 372 -19 378
rect 115 372 173 378
rect 307 372 365 378
rect 499 372 557 378
rect 691 372 749 378
rect 883 372 941 378
rect -845 338 -833 372
rect -653 338 -641 372
rect -461 338 -449 372
rect -269 338 -257 372
rect -77 338 -65 372
rect 115 338 127 372
rect 307 338 319 372
rect 499 338 511 372
rect 691 338 703 372
rect 883 338 895 372
rect -845 332 -787 338
rect -653 332 -595 338
rect -461 332 -403 338
rect -269 332 -211 338
rect -77 332 -19 338
rect 115 332 173 338
rect 307 332 365 338
rect 499 332 557 338
rect 691 332 749 338
rect 883 332 941 338
rect -941 -338 -883 -332
rect -749 -338 -691 -332
rect -557 -338 -499 -332
rect -365 -338 -307 -332
rect -173 -338 -115 -332
rect 19 -338 77 -332
rect 211 -338 269 -332
rect 403 -338 461 -332
rect 595 -338 653 -332
rect 787 -338 845 -332
rect -941 -372 -929 -338
rect -749 -372 -737 -338
rect -557 -372 -545 -338
rect -365 -372 -353 -338
rect -173 -372 -161 -338
rect 19 -372 31 -338
rect 211 -372 223 -338
rect 403 -372 415 -338
rect 595 -372 607 -338
rect 787 -372 799 -338
rect -941 -378 -883 -372
rect -749 -378 -691 -372
rect -557 -378 -499 -372
rect -365 -378 -307 -372
rect -173 -378 -115 -372
rect 19 -378 77 -372
rect 211 -378 269 -372
rect 403 -378 461 -372
rect 595 -378 653 -372
rect 787 -378 845 -372
<< pwell >>
rect -1127 -510 1127 510
<< nmos >>
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
<< ndiff >>
rect -989 288 -927 300
rect -989 -288 -977 288
rect -943 -288 -927 288
rect -989 -300 -927 -288
rect -897 288 -831 300
rect -897 -288 -881 288
rect -847 -288 -831 288
rect -897 -300 -831 -288
rect -801 288 -735 300
rect -801 -288 -785 288
rect -751 -288 -735 288
rect -801 -300 -735 -288
rect -705 288 -639 300
rect -705 -288 -689 288
rect -655 -288 -639 288
rect -705 -300 -639 -288
rect -609 288 -543 300
rect -609 -288 -593 288
rect -559 -288 -543 288
rect -609 -300 -543 -288
rect -513 288 -447 300
rect -513 -288 -497 288
rect -463 -288 -447 288
rect -513 -300 -447 -288
rect -417 288 -351 300
rect -417 -288 -401 288
rect -367 -288 -351 288
rect -417 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 417 300
rect 351 -288 367 288
rect 401 -288 417 288
rect 351 -300 417 -288
rect 447 288 513 300
rect 447 -288 463 288
rect 497 -288 513 288
rect 447 -300 513 -288
rect 543 288 609 300
rect 543 -288 559 288
rect 593 -288 609 288
rect 543 -300 609 -288
rect 639 288 705 300
rect 639 -288 655 288
rect 689 -288 705 288
rect 639 -300 705 -288
rect 735 288 801 300
rect 735 -288 751 288
rect 785 -288 801 288
rect 735 -300 801 -288
rect 831 288 897 300
rect 831 -288 847 288
rect 881 -288 897 288
rect 831 -300 897 -288
rect 927 288 989 300
rect 927 -288 943 288
rect 977 -288 989 288
rect 927 -300 989 -288
<< ndiffc >>
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
<< psubdiff >>
rect -1091 440 -995 474
rect 995 440 1091 474
rect -1091 378 -1057 440
rect 1057 378 1091 440
rect -1091 -440 -1057 -378
rect 1057 -440 1091 -378
rect -1091 -474 -995 -440
rect 995 -474 1091 -440
<< psubdiffcont >>
rect -995 440 995 474
rect -1091 -378 -1057 378
rect 1057 -378 1091 378
rect -995 -474 995 -440
<< poly >>
rect -849 372 -783 388
rect -849 338 -833 372
rect -799 338 -783 372
rect -927 300 -897 326
rect -849 322 -783 338
rect -657 372 -591 388
rect -657 338 -641 372
rect -607 338 -591 372
rect -831 300 -801 322
rect -735 300 -705 326
rect -657 322 -591 338
rect -465 372 -399 388
rect -465 338 -449 372
rect -415 338 -399 372
rect -639 300 -609 322
rect -543 300 -513 326
rect -465 322 -399 338
rect -273 372 -207 388
rect -273 338 -257 372
rect -223 338 -207 372
rect -447 300 -417 322
rect -351 300 -321 326
rect -273 322 -207 338
rect -81 372 -15 388
rect -81 338 -65 372
rect -31 338 -15 372
rect -255 300 -225 322
rect -159 300 -129 326
rect -81 322 -15 338
rect 111 372 177 388
rect 111 338 127 372
rect 161 338 177 372
rect -63 300 -33 322
rect 33 300 63 326
rect 111 322 177 338
rect 303 372 369 388
rect 303 338 319 372
rect 353 338 369 372
rect 129 300 159 322
rect 225 300 255 326
rect 303 322 369 338
rect 495 372 561 388
rect 495 338 511 372
rect 545 338 561 372
rect 321 300 351 322
rect 417 300 447 326
rect 495 322 561 338
rect 687 372 753 388
rect 687 338 703 372
rect 737 338 753 372
rect 513 300 543 322
rect 609 300 639 326
rect 687 322 753 338
rect 879 372 945 388
rect 879 338 895 372
rect 929 338 945 372
rect 705 300 735 322
rect 801 300 831 326
rect 879 322 945 338
rect 897 300 927 322
rect -927 -322 -897 -300
rect -945 -338 -879 -322
rect -831 -326 -801 -300
rect -735 -322 -705 -300
rect -945 -372 -929 -338
rect -895 -372 -879 -338
rect -945 -388 -879 -372
rect -753 -338 -687 -322
rect -639 -326 -609 -300
rect -543 -322 -513 -300
rect -753 -372 -737 -338
rect -703 -372 -687 -338
rect -753 -388 -687 -372
rect -561 -338 -495 -322
rect -447 -326 -417 -300
rect -351 -322 -321 -300
rect -561 -372 -545 -338
rect -511 -372 -495 -338
rect -561 -388 -495 -372
rect -369 -338 -303 -322
rect -255 -326 -225 -300
rect -159 -322 -129 -300
rect -369 -372 -353 -338
rect -319 -372 -303 -338
rect -369 -388 -303 -372
rect -177 -338 -111 -322
rect -63 -326 -33 -300
rect 33 -322 63 -300
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect -177 -388 -111 -372
rect 15 -338 81 -322
rect 129 -326 159 -300
rect 225 -322 255 -300
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 15 -388 81 -372
rect 207 -338 273 -322
rect 321 -326 351 -300
rect 417 -322 447 -300
rect 207 -372 223 -338
rect 257 -372 273 -338
rect 207 -388 273 -372
rect 399 -338 465 -322
rect 513 -326 543 -300
rect 609 -322 639 -300
rect 399 -372 415 -338
rect 449 -372 465 -338
rect 399 -388 465 -372
rect 591 -338 657 -322
rect 705 -326 735 -300
rect 801 -322 831 -300
rect 591 -372 607 -338
rect 641 -372 657 -338
rect 591 -388 657 -372
rect 783 -338 849 -322
rect 897 -326 927 -300
rect 783 -372 799 -338
rect 833 -372 849 -338
rect 783 -388 849 -372
<< polycont >>
rect -833 338 -799 372
rect -641 338 -607 372
rect -449 338 -415 372
rect -257 338 -223 372
rect -65 338 -31 372
rect 127 338 161 372
rect 319 338 353 372
rect 511 338 545 372
rect 703 338 737 372
rect 895 338 929 372
rect -929 -372 -895 -338
rect -737 -372 -703 -338
rect -545 -372 -511 -338
rect -353 -372 -319 -338
rect -161 -372 -127 -338
rect 31 -372 65 -338
rect 223 -372 257 -338
rect 415 -372 449 -338
rect 607 -372 641 -338
rect 799 -372 833 -338
<< locali >>
rect -1091 440 -995 474
rect 995 440 1091 474
rect -1091 378 -1057 440
rect 1057 378 1091 440
rect -849 338 -833 372
rect -799 338 -783 372
rect -657 338 -641 372
rect -607 338 -591 372
rect -465 338 -449 372
rect -415 338 -399 372
rect -273 338 -257 372
rect -223 338 -207 372
rect -81 338 -65 372
rect -31 338 -15 372
rect 111 338 127 372
rect 161 338 177 372
rect 303 338 319 372
rect 353 338 369 372
rect 495 338 511 372
rect 545 338 561 372
rect 687 338 703 372
rect 737 338 753 372
rect 879 338 895 372
rect 929 338 945 372
rect -977 288 -943 304
rect -977 -304 -943 -288
rect -881 288 -847 304
rect -881 -304 -847 -288
rect -785 288 -751 304
rect -785 -304 -751 -288
rect -689 288 -655 304
rect -689 -304 -655 -288
rect -593 288 -559 304
rect -593 -304 -559 -288
rect -497 288 -463 304
rect -497 -304 -463 -288
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect 463 288 497 304
rect 463 -304 497 -288
rect 559 288 593 304
rect 559 -304 593 -288
rect 655 288 689 304
rect 655 -304 689 -288
rect 751 288 785 304
rect 751 -304 785 -288
rect 847 288 881 304
rect 847 -304 881 -288
rect 943 288 977 304
rect 943 -304 977 -288
rect -945 -372 -929 -338
rect -895 -372 -879 -338
rect -753 -372 -737 -338
rect -703 -372 -687 -338
rect -561 -372 -545 -338
rect -511 -372 -495 -338
rect -369 -372 -353 -338
rect -319 -372 -303 -338
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 207 -372 223 -338
rect 257 -372 273 -338
rect 399 -372 415 -338
rect 449 -372 465 -338
rect 591 -372 607 -338
rect 641 -372 657 -338
rect 783 -372 799 -338
rect 833 -372 849 -338
rect -1091 -440 -1057 -378
rect 1057 -440 1091 -378
rect -1091 -474 -995 -440
rect 995 -474 1091 -440
<< viali >>
rect -833 338 -799 372
rect -641 338 -607 372
rect -449 338 -415 372
rect -257 338 -223 372
rect -65 338 -31 372
rect 127 338 161 372
rect 319 338 353 372
rect 511 338 545 372
rect 703 338 737 372
rect 895 338 929 372
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect -929 -372 -895 -338
rect -737 -372 -703 -338
rect -545 -372 -511 -338
rect -353 -372 -319 -338
rect -161 -372 -127 -338
rect 31 -372 65 -338
rect 223 -372 257 -338
rect 415 -372 449 -338
rect 607 -372 641 -338
rect 799 -372 833 -338
<< metal1 >>
rect -845 372 -787 378
rect -845 338 -833 372
rect -799 338 -787 372
rect -845 332 -787 338
rect -653 372 -595 378
rect -653 338 -641 372
rect -607 338 -595 372
rect -653 332 -595 338
rect -461 372 -403 378
rect -461 338 -449 372
rect -415 338 -403 372
rect -461 332 -403 338
rect -269 372 -211 378
rect -269 338 -257 372
rect -223 338 -211 372
rect -269 332 -211 338
rect -77 372 -19 378
rect -77 338 -65 372
rect -31 338 -19 372
rect -77 332 -19 338
rect 115 372 173 378
rect 115 338 127 372
rect 161 338 173 372
rect 115 332 173 338
rect 307 372 365 378
rect 307 338 319 372
rect 353 338 365 372
rect 307 332 365 338
rect 499 372 557 378
rect 499 338 511 372
rect 545 338 557 372
rect 499 332 557 338
rect 691 372 749 378
rect 691 338 703 372
rect 737 338 749 372
rect 691 332 749 338
rect 883 372 941 378
rect 883 338 895 372
rect 929 338 941 372
rect 883 332 941 338
rect -983 288 -937 300
rect -983 -288 -977 288
rect -943 -288 -937 288
rect -983 -300 -937 -288
rect -887 288 -841 300
rect -887 -288 -881 288
rect -847 -288 -841 288
rect -887 -300 -841 -288
rect -791 288 -745 300
rect -791 -288 -785 288
rect -751 -288 -745 288
rect -791 -300 -745 -288
rect -695 288 -649 300
rect -695 -288 -689 288
rect -655 -288 -649 288
rect -695 -300 -649 -288
rect -599 288 -553 300
rect -599 -288 -593 288
rect -559 -288 -553 288
rect -599 -300 -553 -288
rect -503 288 -457 300
rect -503 -288 -497 288
rect -463 -288 -457 288
rect -503 -300 -457 -288
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect 457 288 503 300
rect 457 -288 463 288
rect 497 -288 503 288
rect 457 -300 503 -288
rect 553 288 599 300
rect 553 -288 559 288
rect 593 -288 599 288
rect 553 -300 599 -288
rect 649 288 695 300
rect 649 -288 655 288
rect 689 -288 695 288
rect 649 -300 695 -288
rect 745 288 791 300
rect 745 -288 751 288
rect 785 -288 791 288
rect 745 -300 791 -288
rect 841 288 887 300
rect 841 -288 847 288
rect 881 -288 887 288
rect 841 -300 887 -288
rect 937 288 983 300
rect 937 -288 943 288
rect 977 -288 983 288
rect 937 -300 983 -288
rect -941 -338 -883 -332
rect -941 -372 -929 -338
rect -895 -372 -883 -338
rect -941 -378 -883 -372
rect -749 -338 -691 -332
rect -749 -372 -737 -338
rect -703 -372 -691 -338
rect -749 -378 -691 -372
rect -557 -338 -499 -332
rect -557 -372 -545 -338
rect -511 -372 -499 -338
rect -557 -378 -499 -372
rect -365 -338 -307 -332
rect -365 -372 -353 -338
rect -319 -372 -307 -338
rect -365 -378 -307 -372
rect -173 -338 -115 -332
rect -173 -372 -161 -338
rect -127 -372 -115 -338
rect -173 -378 -115 -372
rect 19 -338 77 -332
rect 19 -372 31 -338
rect 65 -372 77 -338
rect 19 -378 77 -372
rect 211 -338 269 -332
rect 211 -372 223 -338
rect 257 -372 269 -338
rect 211 -378 269 -372
rect 403 -338 461 -332
rect 403 -372 415 -338
rect 449 -372 461 -338
rect 403 -378 461 -372
rect 595 -338 653 -332
rect 595 -372 607 -338
rect 641 -372 653 -338
rect 595 -378 653 -372
rect 787 -338 845 -332
rect 787 -372 799 -338
rect 833 -372 845 -338
rect 787 -378 845 -372
<< properties >>
string FIXED_BBOX -1074 -457 1074 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
