magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -365 372 -307 378
rect -173 372 -115 378
rect 19 372 77 378
rect 211 372 269 378
rect 403 372 461 378
rect -365 338 -353 372
rect -173 338 -161 372
rect 19 338 31 372
rect 211 338 223 372
rect 403 338 415 372
rect -365 332 -307 338
rect -173 332 -115 338
rect 19 332 77 338
rect 211 332 269 338
rect 403 332 461 338
rect -461 -338 -403 -332
rect -269 -338 -211 -332
rect -77 -338 -19 -332
rect 115 -338 173 -332
rect 307 -338 365 -332
rect -461 -372 -449 -338
rect -269 -372 -257 -338
rect -77 -372 -65 -338
rect 115 -372 127 -338
rect 307 -372 319 -338
rect -461 -378 -403 -372
rect -269 -378 -211 -372
rect -77 -378 -19 -372
rect 115 -378 173 -372
rect 307 -378 365 -372
<< pwell >>
rect -647 -510 647 510
<< nmos >>
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
<< ndiff >>
rect -509 288 -447 300
rect -509 -288 -497 288
rect -463 -288 -447 288
rect -509 -300 -447 -288
rect -417 288 -351 300
rect -417 -288 -401 288
rect -367 -288 -351 288
rect -417 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 417 300
rect 351 -288 367 288
rect 401 -288 417 288
rect 351 -300 417 -288
rect 447 288 509 300
rect 447 -288 463 288
rect 497 -288 509 288
rect 447 -300 509 -288
<< ndiffc >>
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
<< psubdiff >>
rect -611 440 -515 474
rect 515 440 611 474
rect -611 378 -577 440
rect 577 378 611 440
rect -611 -440 -577 -378
rect 577 -440 611 -378
rect -611 -474 -515 -440
rect 515 -474 611 -440
<< psubdiffcont >>
rect -515 440 515 474
rect -611 -378 -577 378
rect 577 -378 611 378
rect -515 -474 515 -440
<< poly >>
rect -369 372 -303 388
rect -369 338 -353 372
rect -319 338 -303 372
rect -447 300 -417 326
rect -369 322 -303 338
rect -177 372 -111 388
rect -177 338 -161 372
rect -127 338 -111 372
rect -351 300 -321 322
rect -255 300 -225 326
rect -177 322 -111 338
rect 15 372 81 388
rect 15 338 31 372
rect 65 338 81 372
rect -159 300 -129 322
rect -63 300 -33 326
rect 15 322 81 338
rect 207 372 273 388
rect 207 338 223 372
rect 257 338 273 372
rect 33 300 63 322
rect 129 300 159 326
rect 207 322 273 338
rect 399 372 465 388
rect 399 338 415 372
rect 449 338 465 372
rect 225 300 255 322
rect 321 300 351 326
rect 399 322 465 338
rect 417 300 447 322
rect -447 -322 -417 -300
rect -465 -338 -399 -322
rect -351 -326 -321 -300
rect -255 -322 -225 -300
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -465 -388 -399 -372
rect -273 -338 -207 -322
rect -159 -326 -129 -300
rect -63 -322 -33 -300
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -273 -388 -207 -372
rect -81 -338 -15 -322
rect 33 -326 63 -300
rect 129 -322 159 -300
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect -81 -388 -15 -372
rect 111 -338 177 -322
rect 225 -326 255 -300
rect 321 -322 351 -300
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 111 -388 177 -372
rect 303 -338 369 -322
rect 417 -326 447 -300
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 303 -388 369 -372
<< polycont >>
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
<< locali >>
rect -611 440 -515 474
rect 515 440 611 474
rect -611 378 -577 440
rect 577 378 611 440
rect -369 338 -353 372
rect -319 338 -303 372
rect -177 338 -161 372
rect -127 338 -111 372
rect 15 338 31 372
rect 65 338 81 372
rect 207 338 223 372
rect 257 338 273 372
rect 399 338 415 372
rect 449 338 465 372
rect -497 288 -463 304
rect -497 -304 -463 -288
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect 463 288 497 304
rect 463 -304 497 -288
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 303 -372 319 -338
rect 353 -372 369 -338
rect -611 -440 -577 -378
rect 577 -440 611 -378
rect -611 -474 -515 -440
rect 515 -474 611 -440
<< viali >>
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
<< metal1 >>
rect -365 372 -307 378
rect -365 338 -353 372
rect -319 338 -307 372
rect -365 332 -307 338
rect -173 372 -115 378
rect -173 338 -161 372
rect -127 338 -115 372
rect -173 332 -115 338
rect 19 372 77 378
rect 19 338 31 372
rect 65 338 77 372
rect 19 332 77 338
rect 211 372 269 378
rect 211 338 223 372
rect 257 338 269 372
rect 211 332 269 338
rect 403 372 461 378
rect 403 338 415 372
rect 449 338 461 372
rect 403 332 461 338
rect -503 288 -457 300
rect -503 -288 -497 288
rect -463 -288 -457 288
rect -503 -300 -457 -288
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect 457 288 503 300
rect 457 -288 463 288
rect 497 -288 503 288
rect 457 -300 503 -288
rect -461 -338 -403 -332
rect -461 -372 -449 -338
rect -415 -372 -403 -338
rect -461 -378 -403 -372
rect -269 -338 -211 -332
rect -269 -372 -257 -338
rect -223 -372 -211 -338
rect -269 -378 -211 -372
rect -77 -338 -19 -332
rect -77 -372 -65 -338
rect -31 -372 -19 -338
rect -77 -378 -19 -372
rect 115 -338 173 -332
rect 115 -372 127 -338
rect 161 -372 173 -338
rect 115 -378 173 -372
rect 307 -338 365 -332
rect 307 -372 319 -338
rect 353 -372 365 -338
rect 307 -378 365 -372
<< properties >>
string FIXED_BBOX -594 -457 594 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
