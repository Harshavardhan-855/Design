magic
tech sky130A
magscale 1 2
timestamp 1708427081
<< checkpaint >>
rect -1260 17387 16048 19987
rect -1734 11963 16048 17387
rect -2558 -660 16048 11963
rect -2558 -3260 15612 -660
rect -2558 -8684 14750 -3260
<< error_s >>
rect 862 9720 2274 9724
rect 834 9692 2246 9696
rect 931 9631 1029 9651
rect 1079 9631 1113 9653
rect 1237 9631 1316 9659
rect 1320 9655 1322 9669
rect 1623 9655 1626 9669
rect 1320 9651 1392 9655
rect 1414 9651 1500 9655
rect 1320 9637 1511 9651
rect 1513 9637 1626 9655
rect 1760 9649 1802 9655
rect 1750 9647 1802 9649
rect 1653 9637 1720 9647
rect 1749 9637 1802 9647
rect 1092 9627 1107 9631
rect 896 9613 926 9627
rect 1081 9623 1107 9627
rect 931 9613 1029 9617
rect 896 9601 1029 9613
rect 897 9599 1029 9601
rect 1065 9601 1107 9623
rect 1065 9599 1109 9601
rect 902 9597 1029 9599
rect 902 9583 1004 9597
rect 1039 9589 1055 9599
rect 1065 9593 1103 9599
rect 1093 9589 1097 9593
rect 1049 9587 1055 9589
rect 941 9579 971 9583
rect 902 9549 914 9579
rect 936 9572 971 9579
rect 926 9542 971 9572
rect 926 9532 938 9542
rect 950 9535 970 9542
rect 950 9532 978 9535
rect 926 9520 978 9532
rect 847 9517 978 9520
rect 884 9423 896 9489
rect 950 9477 970 9517
rect 984 9460 1004 9583
rect 1041 9561 1067 9587
rect 1025 9460 1030 9539
rect 980 9444 1030 9460
rect 1025 9443 1030 9444
rect 1041 9535 1055 9561
rect 1099 9539 1103 9593
rect 1133 9557 1137 9631
rect 1184 9581 1198 9631
rect 1320 9627 1322 9637
rect 1350 9631 1426 9637
rect 1447 9631 1511 9637
rect 1512 9627 1513 9637
rect 1271 9601 1316 9625
rect 1362 9601 1364 9627
rect 1384 9601 1426 9617
rect 1476 9615 1477 9617
rect 1443 9601 1477 9615
rect 1554 9601 1555 9627
rect 1623 9601 1626 9637
rect 1849 9631 1961 9659
rect 2001 9637 2016 9655
rect 2022 9649 2088 9655
rect 2106 9653 2136 9655
rect 2091 9649 2136 9653
rect 2142 9649 2186 9655
rect 2022 9637 2186 9649
rect 2022 9631 2182 9637
rect 2216 9631 2246 9665
rect 2250 9659 2280 9699
rect 1271 9597 1477 9601
rect 1218 9581 1232 9597
rect 1308 9593 1477 9597
rect 1308 9589 1465 9593
rect 1308 9586 1337 9589
rect 1041 9454 1077 9535
rect 1156 9534 1284 9581
rect 1308 9535 1322 9586
rect 1384 9555 1465 9589
rect 1392 9545 1434 9555
rect 1203 9529 1284 9534
rect 1305 9529 1358 9535
rect 1203 9517 1278 9529
rect 1308 9517 1325 9529
rect 1392 9517 1470 9518
rect 1203 9500 1224 9517
rect 1041 9448 1055 9454
rect 1059 9448 1064 9454
rect 1041 9433 1070 9448
rect 1097 9433 1099 9471
rect 1093 9423 1099 9433
rect 1131 9423 1133 9437
rect 1305 9435 1324 9495
rect 1339 9443 1358 9501
rect 1476 9453 1477 9589
rect 1500 9586 1528 9601
rect 1500 9532 1513 9586
rect 1586 9563 1641 9601
rect 1649 9563 1651 9589
rect 1697 9578 1749 9593
rect 1623 9555 1641 9563
rect 1697 9555 1714 9578
rect 1617 9532 1714 9555
rect 1500 9517 1528 9532
rect 1608 9529 1714 9532
rect 1608 9521 1641 9529
rect 1510 9503 1511 9517
rect 1500 9487 1513 9503
rect 1500 9473 1548 9487
rect 1554 9473 1555 9517
rect 1583 9495 1670 9521
rect 1511 9469 1548 9473
rect 1511 9461 1556 9469
rect 1582 9461 1636 9487
rect 1542 9453 1556 9461
rect 1237 9423 1266 9435
rect 1271 9423 1305 9435
rect 1339 9423 1360 9443
rect 1477 9427 1556 9453
rect 1582 9427 1602 9453
rect 1542 9423 1556 9427
rect 1589 9423 1602 9427
rect 1623 9423 1636 9427
rect 1637 9423 1638 9495
rect 1720 9480 1749 9578
rect 1849 9563 1852 9631
rect 1865 9627 1880 9631
rect 1865 9625 1891 9627
rect 1947 9625 1968 9627
rect 1865 9601 1968 9625
rect 2022 9601 2028 9631
rect 2046 9605 2052 9627
rect 2056 9601 2148 9615
rect 2156 9601 2182 9631
rect 1883 9597 1961 9601
rect 1883 9563 1886 9597
rect 1917 9553 1918 9597
rect 2001 9586 2028 9601
rect 2051 9589 2198 9601
rect 2016 9557 2028 9586
rect 2056 9557 2062 9589
rect 2073 9586 2198 9589
rect 2016 9554 2022 9557
rect 2088 9555 2182 9586
rect 1750 9538 1883 9545
rect 1917 9538 1938 9553
rect 2010 9545 2062 9554
rect 1750 9529 1938 9538
rect 1841 9522 1846 9529
rect 1768 9511 1849 9522
rect 1876 9511 1938 9529
rect 1997 9523 2062 9545
rect 2088 9539 2122 9555
rect 2136 9539 2142 9555
rect 1750 9508 1938 9511
rect 1750 9495 1883 9508
rect 1705 9474 1749 9480
rect 1768 9475 1849 9495
rect 1697 9467 1800 9474
rect 1805 9467 1849 9475
rect 1955 9467 1971 9477
rect 1697 9465 1993 9467
rect 1723 9462 1993 9465
rect 1997 9462 2005 9511
rect 2016 9510 2022 9523
rect 2044 9510 2062 9520
rect 2101 9510 2122 9539
rect 2156 9521 2182 9555
rect 2135 9510 2156 9521
rect 2012 9484 2156 9510
rect 2186 9487 2198 9586
rect 2284 9583 2341 9607
rect 2397 9583 2460 9607
rect 2521 9585 2573 9607
rect 2593 9594 2620 9607
rect 2593 9585 2635 9594
rect 2250 9549 2341 9573
rect 2376 9539 2385 9558
rect 2397 9539 2426 9573
rect 2592 9553 2599 9583
rect 2620 9579 2635 9585
rect 2660 9583 2761 9597
rect 2834 9583 2836 9617
rect 2620 9553 2646 9579
rect 2701 9563 2731 9579
rect 2868 9569 2870 9633
rect 3698 9624 5110 9628
rect 3670 9596 5082 9600
rect 2558 9538 2599 9553
rect 2169 9484 2198 9487
rect 2012 9463 2198 9484
rect 2031 9462 2039 9463
rect 821 9419 896 9423
rect 903 9419 1192 9423
rect 821 9409 1192 9419
rect 821 9385 896 9409
rect 903 9385 1192 9409
rect 1237 9411 1428 9423
rect 1451 9411 1561 9423
rect 1589 9419 1708 9423
rect 1237 9403 1561 9411
rect 821 9381 1192 9385
rect 1242 9381 1561 9403
rect 1591 9403 1708 9419
rect 1723 9403 2044 9462
rect 1591 9401 2044 9403
rect 2052 9445 2198 9463
rect 2345 9496 2401 9511
rect 2431 9505 2460 9515
rect 2541 9511 2549 9520
rect 2052 9423 2122 9445
rect 2135 9437 2198 9445
rect 2135 9423 2156 9437
rect 2169 9423 2198 9437
rect 2203 9423 2224 9453
rect 2283 9431 2343 9443
rect 2345 9442 2380 9496
rect 2385 9442 2401 9496
rect 2495 9489 2549 9511
rect 2573 9489 2599 9538
rect 2626 9489 2633 9553
rect 2694 9551 2761 9563
rect 2670 9549 2761 9551
rect 2670 9521 2697 9549
rect 2701 9541 2744 9549
rect 2762 9541 2792 9551
rect 2701 9521 2731 9541
rect 2761 9529 2792 9541
rect 2670 9489 2700 9521
rect 2762 9489 2792 9529
rect 2847 9521 2930 9553
rect 2345 9431 2401 9442
rect 2345 9427 2358 9431
rect 2370 9427 2401 9431
rect 2425 9423 2431 9483
rect 2495 9473 2599 9489
rect 2532 9439 2599 9473
rect 2491 9423 2494 9439
rect 2532 9427 2593 9439
rect 2623 9427 2701 9489
rect 2731 9439 2792 9489
rect 2797 9473 2807 9507
rect 2892 9499 2912 9501
rect 2943 9499 2946 9535
rect 2953 9521 3022 9553
rect 3091 9535 3222 9563
rect 3255 9547 3477 9559
rect 3315 9535 3477 9547
rect 2844 9469 2854 9473
rect 2858 9469 2878 9489
rect 2892 9469 2953 9499
rect 2807 9439 2953 9469
rect 2731 9427 2953 9439
rect 2977 9444 2980 9521
rect 3125 9501 3188 9529
rect 3396 9525 3417 9531
rect 2977 9435 3043 9444
rect 2532 9423 3048 9427
rect 2052 9413 2535 9423
rect 2052 9401 2094 9413
rect 1567 9381 1582 9397
rect 1591 9381 2010 9401
rect 2022 9399 2049 9401
rect 2020 9381 2049 9399
rect 2101 9381 2535 9413
rect 2573 9381 3048 9423
rect 821 9371 3048 9381
rect 3091 9403 3111 9501
rect 3125 9403 3145 9501
rect 3252 9490 3270 9505
rect 3315 9501 3443 9525
rect 3495 9505 3525 9531
rect 3585 9501 3591 9525
rect 3620 9505 3631 9546
rect 3767 9535 3865 9555
rect 3915 9535 3949 9557
rect 4073 9535 4152 9563
rect 4156 9559 4158 9573
rect 4459 9559 4462 9573
rect 4156 9555 4228 9559
rect 4250 9555 4336 9559
rect 4156 9541 4347 9555
rect 4349 9541 4462 9559
rect 4596 9553 4638 9559
rect 4586 9551 4638 9553
rect 4489 9541 4556 9551
rect 4585 9541 4638 9551
rect 3334 9490 3354 9501
rect 3427 9491 3447 9501
rect 3252 9475 3255 9490
rect 3244 9472 3294 9475
rect 3334 9472 3339 9490
rect 3375 9472 3378 9491
rect 3409 9472 3412 9491
rect 3437 9473 3447 9491
rect 3551 9473 3557 9501
rect 3585 9491 3619 9501
rect 3585 9475 3591 9491
rect 3638 9475 3643 9535
rect 3426 9472 3447 9473
rect 3244 9443 3467 9472
rect 3252 9441 3265 9443
rect 3210 9436 3265 9441
rect 3278 9441 3467 9443
rect 3525 9441 3557 9473
rect 3672 9449 3677 9535
rect 3928 9531 3943 9535
rect 3732 9517 3762 9531
rect 3917 9527 3943 9531
rect 3767 9517 3865 9521
rect 3732 9505 3865 9517
rect 3733 9503 3865 9505
rect 3901 9505 3943 9527
rect 3901 9503 3945 9505
rect 3738 9501 3865 9503
rect 3738 9487 3840 9501
rect 3875 9493 3891 9503
rect 3901 9497 3939 9503
rect 3929 9493 3933 9497
rect 3885 9491 3891 9493
rect 3777 9483 3807 9487
rect 3738 9453 3750 9483
rect 3772 9476 3807 9483
rect 3762 9446 3807 9476
rect 3210 9421 3270 9436
rect 3278 9425 3495 9441
rect 3525 9436 3555 9441
rect 3762 9436 3774 9446
rect 3786 9439 3806 9446
rect 3786 9436 3814 9439
rect 3309 9421 3406 9425
rect 3409 9421 3412 9425
rect 3426 9421 3495 9425
rect 3501 9421 3523 9435
rect 3525 9421 3570 9436
rect 3762 9424 3814 9436
rect 3683 9421 3814 9424
rect 3210 9409 3263 9421
rect 3297 9409 3699 9421
rect 3249 9403 3263 9409
rect 3283 9403 3699 9409
rect 821 9365 3090 9371
rect 941 9355 968 9365
rect 981 9355 1013 9365
rect 1025 9355 1030 9365
rect 1059 9355 1064 9365
rect 889 9351 941 9355
rect 971 9351 1064 9355
rect 889 9341 1025 9351
rect 889 9317 967 9341
rect 971 9340 1025 9341
rect 981 9317 1025 9340
rect 1059 9343 1064 9351
rect 889 9305 1031 9317
rect 889 9279 991 9305
rect 871 9275 991 9279
rect 828 9271 991 9275
rect 828 9257 993 9271
rect 941 9245 957 9257
rect 965 9245 993 9257
rect 965 9241 991 9245
rect 1007 9241 1031 9305
rect 1059 9271 1065 9343
rect 1097 9293 1099 9365
rect 1101 9271 1107 9333
rect 1131 9275 1133 9365
rect 1277 9355 1310 9365
rect 1177 9353 1307 9355
rect 1177 9340 1192 9353
rect 1197 9343 1307 9353
rect 1213 9341 1307 9343
rect 1139 9275 1145 9295
rect 1175 9286 1211 9333
rect 1225 9309 1307 9341
rect 1311 9319 1339 9365
rect 1567 9355 1582 9365
rect 1601 9355 1636 9363
rect 1341 9343 1360 9355
rect 1519 9345 1636 9355
rect 1501 9343 1636 9345
rect 1670 9355 1768 9365
rect 1791 9355 1841 9365
rect 1670 9343 1841 9355
rect 1341 9328 1471 9343
rect 1341 9317 1451 9328
rect 1225 9293 1279 9309
rect 1345 9297 1375 9317
rect 1225 9289 1255 9293
rect 1321 9289 1375 9297
rect 1379 9311 1451 9317
rect 1465 9311 1471 9328
rect 1475 9340 1616 9343
rect 1693 9340 1709 9343
rect 1475 9311 1547 9340
rect 1379 9289 1519 9311
rect 1561 9289 1591 9340
rect 1601 9289 1616 9340
rect 1708 9303 1709 9340
rect 1718 9319 1841 9343
rect 1739 9303 1841 9319
rect 1749 9289 1779 9303
rect 1225 9286 1794 9289
rect 1041 9241 1065 9271
rect 1131 9245 1171 9275
rect 1175 9271 1794 9286
rect 1831 9275 1836 9303
rect 1865 9279 1870 9365
rect 1871 9343 1937 9365
rect 2010 9343 2012 9365
rect 2101 9355 2122 9365
rect 2135 9355 2175 9365
rect 2203 9363 2224 9365
rect 2095 9353 2156 9355
rect 1871 9303 1940 9343
rect 1995 9331 2054 9343
rect 2079 9331 2156 9353
rect 1995 9328 2136 9331
rect 2010 9319 2136 9328
rect 2010 9303 2049 9319
rect 2079 9303 2136 9319
rect 1871 9281 1876 9303
rect 1938 9281 1940 9303
rect 1885 9279 1919 9281
rect 1979 9275 2088 9303
rect 2106 9281 2136 9303
rect 2169 9281 2190 9309
rect 1237 9245 1277 9271
rect 1280 9245 1297 9271
rect 1321 9267 1352 9271
rect 1379 9267 1485 9271
rect 1321 9245 1351 9267
rect 1375 9251 1485 9267
rect 1519 9257 1553 9271
rect 1601 9251 1616 9271
rect 1375 9245 1451 9251
rect 1749 9247 1779 9271
rect 1823 9247 1836 9275
rect 2106 9271 2121 9281
rect 1379 9243 1451 9245
rect 1723 9245 1789 9247
rect 1841 9245 1846 9271
rect 1968 9245 1970 9271
rect 2052 9269 2079 9271
rect 1723 9241 1755 9245
rect 1757 9241 1789 9245
rect 1978 9241 2012 9269
rect 2046 9241 2088 9269
rect 2145 9245 2190 9281
rect 2169 9241 2190 9245
rect 2203 9241 2224 9324
rect 2246 9317 3090 9365
rect 3091 9357 3699 9403
rect 3101 9335 3699 9357
rect 2322 9305 2432 9317
rect 2344 9286 2432 9305
rect 2329 9275 2446 9286
rect 2451 9283 2459 9317
rect 2463 9305 2467 9317
rect 2301 9271 2446 9275
rect 2485 9275 2493 9317
rect 2521 9305 2670 9317
rect 2501 9275 2505 9305
rect 2521 9293 2579 9305
rect 2521 9287 2573 9293
rect 2585 9287 2670 9305
rect 2677 9287 2694 9317
rect 2700 9287 2731 9317
rect 2836 9287 3090 9317
rect 2521 9282 3090 9287
rect 3143 9327 3699 9335
rect 3720 9327 3732 9393
rect 3786 9381 3806 9421
rect 3820 9364 3840 9487
rect 3877 9465 3903 9491
rect 3861 9364 3866 9443
rect 3816 9348 3866 9364
rect 3861 9347 3866 9348
rect 3877 9439 3891 9465
rect 3935 9443 3939 9497
rect 3969 9461 3973 9535
rect 4020 9485 4034 9535
rect 4156 9531 4158 9541
rect 4186 9535 4262 9541
rect 4283 9535 4347 9541
rect 4348 9531 4349 9541
rect 4107 9505 4152 9529
rect 4198 9505 4200 9531
rect 4220 9505 4262 9521
rect 4312 9519 4313 9521
rect 4279 9505 4313 9519
rect 4390 9505 4391 9531
rect 4459 9505 4462 9541
rect 4685 9535 4797 9563
rect 4837 9541 4852 9559
rect 4858 9553 4924 9559
rect 4942 9557 4972 9559
rect 4927 9553 4972 9557
rect 4978 9553 5022 9559
rect 4858 9541 5022 9553
rect 4858 9535 5018 9541
rect 5052 9535 5082 9569
rect 5086 9563 5116 9603
rect 4107 9501 4313 9505
rect 4054 9485 4068 9501
rect 4144 9497 4313 9501
rect 4144 9493 4301 9497
rect 4144 9490 4173 9493
rect 3877 9358 3913 9439
rect 3992 9438 4120 9485
rect 4144 9439 4158 9490
rect 4220 9459 4301 9493
rect 4228 9449 4270 9459
rect 4039 9433 4120 9438
rect 4141 9433 4194 9439
rect 4039 9421 4114 9433
rect 4144 9421 4161 9433
rect 4228 9421 4306 9422
rect 4039 9404 4060 9421
rect 3877 9352 3891 9358
rect 3895 9352 3900 9358
rect 3877 9337 3906 9352
rect 3933 9337 3935 9375
rect 3929 9327 3935 9337
rect 3967 9327 3969 9341
rect 4141 9339 4160 9399
rect 4175 9347 4194 9405
rect 4312 9357 4313 9493
rect 4336 9490 4364 9505
rect 4336 9436 4349 9490
rect 4422 9467 4477 9505
rect 4485 9467 4487 9493
rect 4533 9482 4585 9497
rect 4459 9459 4477 9467
rect 4533 9459 4550 9482
rect 4453 9436 4550 9459
rect 4336 9421 4364 9436
rect 4444 9433 4550 9436
rect 4444 9425 4477 9433
rect 4346 9407 4347 9421
rect 4336 9391 4349 9407
rect 4336 9377 4384 9391
rect 4390 9377 4391 9421
rect 4419 9399 4506 9425
rect 4347 9373 4384 9377
rect 4347 9365 4392 9373
rect 4418 9365 4472 9391
rect 4378 9357 4392 9365
rect 4073 9327 4102 9339
rect 4107 9327 4141 9339
rect 4175 9327 4196 9347
rect 4313 9331 4392 9357
rect 4418 9331 4438 9357
rect 4378 9327 4392 9331
rect 4425 9327 4438 9331
rect 4459 9327 4472 9331
rect 4473 9327 4474 9399
rect 4556 9384 4585 9482
rect 4685 9467 4688 9535
rect 4701 9531 4716 9535
rect 4701 9529 4727 9531
rect 4783 9529 4804 9531
rect 4701 9505 4804 9529
rect 4858 9505 4864 9535
rect 4882 9509 4888 9531
rect 4892 9505 4984 9519
rect 4992 9505 5018 9535
rect 5409 9511 5439 9525
rect 4719 9501 4797 9505
rect 4719 9467 4722 9501
rect 4753 9457 4754 9501
rect 4837 9490 4864 9505
rect 4887 9493 5034 9505
rect 4852 9461 4864 9490
rect 4892 9461 4898 9493
rect 4909 9490 5034 9493
rect 4852 9458 4858 9461
rect 4924 9459 5018 9490
rect 4586 9442 4719 9449
rect 4753 9442 4774 9457
rect 4846 9449 4898 9458
rect 4586 9433 4774 9442
rect 4677 9426 4682 9433
rect 4604 9415 4685 9426
rect 4712 9415 4774 9433
rect 4833 9427 4898 9449
rect 4924 9443 4958 9459
rect 4972 9443 4978 9459
rect 4586 9412 4774 9415
rect 4586 9399 4719 9412
rect 4541 9378 4585 9384
rect 4604 9379 4685 9399
rect 4533 9371 4636 9378
rect 4641 9371 4685 9379
rect 4791 9371 4807 9381
rect 4533 9369 4829 9371
rect 4559 9366 4829 9369
rect 4833 9366 4841 9415
rect 4852 9414 4858 9427
rect 4880 9414 4898 9424
rect 4937 9414 4958 9443
rect 4992 9425 5018 9459
rect 4971 9414 4992 9425
rect 4848 9388 4992 9414
rect 5022 9391 5034 9490
rect 5120 9487 5146 9511
rect 5199 9487 5296 9511
rect 5357 9489 5456 9511
rect 5251 9483 5256 9487
rect 5086 9453 5146 9477
rect 5199 9457 5267 9477
rect 5293 9457 5298 9483
rect 5005 9388 5034 9391
rect 4848 9367 5034 9388
rect 4867 9366 4875 9367
rect 3143 9323 3732 9327
rect 3739 9323 4028 9327
rect 3143 9313 4028 9323
rect 3143 9289 3732 9313
rect 3739 9289 4028 9313
rect 4073 9315 4264 9327
rect 4287 9315 4397 9327
rect 4425 9323 4544 9327
rect 4073 9307 4397 9315
rect 3143 9285 4028 9289
rect 4078 9285 4397 9307
rect 4427 9307 4544 9323
rect 4559 9307 4880 9366
rect 4427 9305 4880 9307
rect 4888 9349 5034 9367
rect 5157 9442 5175 9457
rect 5187 9453 5293 9457
rect 5187 9442 5209 9453
rect 5157 9416 5160 9442
rect 5202 9427 5209 9442
rect 5212 9443 5293 9453
rect 5212 9441 5228 9443
rect 5230 9442 5271 9443
rect 5230 9441 5261 9442
rect 5157 9385 5165 9416
rect 4888 9327 4958 9349
rect 4971 9341 5034 9349
rect 4971 9327 4992 9341
rect 5005 9327 5034 9341
rect 5039 9327 5060 9357
rect 5157 9343 5179 9385
rect 5199 9343 5227 9409
rect 5157 9335 5227 9343
rect 5146 9327 5179 9335
rect 4888 9317 5198 9327
rect 4888 9305 4930 9317
rect 4403 9285 4418 9301
rect 4427 9285 4846 9305
rect 4858 9303 4885 9305
rect 4856 9285 4885 9303
rect 4937 9285 5198 9317
rect 5199 9285 5227 9335
rect 5233 9285 5261 9441
rect 5299 9393 5330 9487
rect 5333 9424 5364 9487
rect 5409 9457 5439 9489
rect 5543 9487 5580 9501
rect 5467 9483 5496 9487
rect 5461 9457 5496 9483
rect 5407 9445 5454 9457
rect 5407 9442 5451 9445
rect 5409 9424 5439 9442
rect 5333 9411 5451 9424
rect 5331 9393 5459 9411
rect 5467 9393 5496 9457
rect 5501 9457 5530 9487
rect 5501 9455 5533 9457
rect 5501 9408 5536 9455
rect 5543 9453 5597 9467
rect 5546 9433 5569 9453
rect 5501 9395 5543 9408
rect 5506 9393 5543 9395
rect 5331 9377 5461 9393
rect 5299 9327 5330 9343
rect 5333 9339 5364 9343
rect 5333 9327 5367 9339
rect 5368 9327 5377 9377
rect 5378 9343 5461 9377
rect 5467 9373 5543 9393
rect 5467 9361 5618 9373
rect 5407 9331 5461 9343
rect 5491 9331 5618 9361
rect 5906 9341 5926 9373
rect 5407 9327 5618 9331
rect 5365 9293 5401 9305
rect 5409 9285 5618 9327
rect 2521 9275 3048 9282
rect 2485 9271 3048 9275
rect 2344 9255 2366 9271
rect 2573 9259 2613 9271
rect 2573 9255 2593 9259
rect 2643 9241 2660 9271
rect 2677 9241 2694 9271
rect 2701 9245 2731 9255
rect 2762 9245 2773 9271
rect 2836 9269 3048 9271
rect 2896 9245 2918 9269
rect 2946 9241 2962 9269
rect 2980 9263 3002 9269
rect 2980 9260 3030 9263
rect 2980 9241 3041 9260
rect 3077 9252 3104 9275
rect 3143 9269 5618 9285
rect 3205 9268 3225 9269
rect 3255 9268 3309 9269
rect 3292 9266 3309 9268
rect 3277 9252 3309 9266
rect 3322 9252 3339 9269
rect 3387 9257 3421 9269
rect 3441 9257 3525 9269
rect 3777 9259 3804 9269
rect 3817 9259 3849 9269
rect 3861 9259 3866 9269
rect 3895 9259 3900 9269
rect 3387 9252 3455 9257
rect 3725 9255 3777 9259
rect 3807 9255 3900 9259
rect 862 9223 991 9241
rect 1097 9227 1171 9241
rect 891 9219 925 9223
rect 1093 9211 1171 9227
rect 1237 9235 1311 9241
rect 1237 9230 1321 9235
rect 1237 9211 1311 9230
rect 1093 9207 1145 9211
rect 1345 9209 1451 9241
rect 1500 9231 1516 9235
rect 1535 9231 1569 9241
rect 1485 9207 1601 9231
rect 1622 9230 1643 9235
rect 1697 9230 1749 9235
rect 1755 9213 1757 9241
rect 1823 9213 1870 9241
rect 2271 9237 2581 9241
rect 2558 9230 2593 9233
rect 2655 9230 2701 9233
rect 2747 9230 2807 9233
rect 2996 9229 3041 9241
rect 3007 9207 3041 9229
rect 3043 9207 3070 9241
rect 3077 9232 3351 9252
rect 3387 9249 3688 9252
rect 3365 9232 3688 9249
rect 3725 9245 3861 9255
rect 1093 9180 1111 9193
rect 1485 9180 1601 9197
rect 862 9176 2274 9180
rect 1093 9173 1111 9176
rect 1485 9173 1601 9176
rect 3077 9173 3104 9232
rect 3292 9225 3297 9232
rect 3322 9227 3339 9232
rect 3365 9231 3551 9232
rect 3363 9229 3551 9231
rect 3365 9227 3551 9229
rect 3364 9225 3548 9227
rect 3365 9224 3548 9225
rect 3560 9224 3585 9232
rect 3108 9204 3351 9224
rect 3365 9223 3660 9224
rect 3407 9211 3660 9223
rect 3408 9204 3660 9211
rect 3725 9221 3803 9245
rect 3807 9244 3861 9245
rect 3817 9221 3861 9244
rect 3895 9247 3900 9255
rect 3725 9209 3867 9221
rect 3408 9193 3421 9204
rect 3460 9197 3526 9204
rect 3489 9193 3526 9197
rect 3560 9193 3585 9204
rect 3325 9191 3355 9193
rect 3597 9159 3631 9193
rect 3635 9179 3669 9195
rect 3725 9183 3827 9209
rect 3707 9179 3827 9183
rect 3635 9175 3827 9179
rect 3635 9161 3829 9175
rect 834 9148 2246 9152
rect 3777 9149 3793 9161
rect 3801 9149 3829 9161
rect 3801 9145 3827 9149
rect 3843 9145 3867 9209
rect 3895 9175 3901 9247
rect 3933 9197 3935 9269
rect 3937 9175 3943 9237
rect 3967 9179 3969 9269
rect 4113 9259 4146 9269
rect 4013 9257 4143 9259
rect 4013 9244 4028 9257
rect 4033 9247 4143 9257
rect 4049 9245 4143 9247
rect 3975 9179 3981 9199
rect 4011 9190 4047 9237
rect 4061 9213 4143 9245
rect 4147 9223 4175 9269
rect 4403 9259 4418 9269
rect 4437 9259 4472 9267
rect 4177 9247 4196 9259
rect 4355 9249 4472 9259
rect 4337 9247 4472 9249
rect 4506 9259 4604 9269
rect 4627 9259 4677 9269
rect 4506 9247 4677 9259
rect 4177 9232 4307 9247
rect 4177 9221 4287 9232
rect 4061 9197 4115 9213
rect 4181 9201 4211 9221
rect 4061 9193 4091 9197
rect 4157 9193 4211 9201
rect 4215 9215 4287 9221
rect 4301 9215 4307 9232
rect 4311 9244 4452 9247
rect 4529 9244 4545 9247
rect 4311 9215 4383 9244
rect 4215 9193 4355 9215
rect 4397 9193 4427 9244
rect 4437 9193 4452 9244
rect 4544 9207 4545 9244
rect 4554 9223 4677 9247
rect 4575 9207 4677 9223
rect 4585 9193 4615 9207
rect 4061 9190 4630 9193
rect 3877 9145 3901 9175
rect 3967 9149 4007 9179
rect 4011 9175 4630 9190
rect 4667 9179 4672 9207
rect 4701 9183 4706 9269
rect 4707 9247 4773 9269
rect 4846 9247 4848 9269
rect 4937 9259 4958 9269
rect 4971 9259 5011 9269
rect 5039 9267 5060 9269
rect 4931 9257 4992 9259
rect 4707 9207 4776 9247
rect 4831 9235 4890 9247
rect 4915 9235 4992 9257
rect 4831 9232 4972 9235
rect 4846 9223 4972 9232
rect 4846 9207 4885 9223
rect 4915 9207 4972 9223
rect 4707 9185 4712 9207
rect 4774 9185 4776 9207
rect 4721 9183 4755 9185
rect 4815 9179 4924 9207
rect 4942 9185 4972 9207
rect 5005 9185 5026 9213
rect 4073 9149 4113 9175
rect 4116 9149 4133 9175
rect 4157 9171 4188 9175
rect 4215 9171 4321 9175
rect 4157 9149 4187 9171
rect 4211 9155 4321 9171
rect 4355 9161 4389 9175
rect 4437 9155 4452 9175
rect 4211 9149 4287 9155
rect 4585 9151 4615 9175
rect 4659 9151 4672 9179
rect 4942 9175 4957 9185
rect 4215 9147 4287 9149
rect 4559 9149 4625 9151
rect 4677 9149 4682 9175
rect 4804 9149 4806 9175
rect 4888 9173 4915 9175
rect 4559 9145 4591 9149
rect 4593 9145 4625 9149
rect 4814 9145 4848 9173
rect 4882 9145 4924 9173
rect 4981 9149 5026 9185
rect 5005 9145 5026 9149
rect 5039 9145 5060 9228
rect 5082 9221 5618 9269
rect 5119 9209 5303 9221
rect 5157 9191 5229 9209
rect 5249 9191 5303 9209
rect 5103 9179 5303 9191
rect 5357 9209 5496 9221
rect 5357 9191 5409 9209
rect 5417 9191 5496 9209
rect 5501 9191 5530 9221
rect 5357 9179 5597 9191
rect 5103 9175 5597 9179
rect 5467 9159 5496 9175
rect 5409 9149 5439 9159
rect 5461 9149 5496 9159
rect 5467 9145 5496 9149
rect 5501 9149 5533 9175
rect 5501 9145 5530 9149
rect 3698 9127 3827 9145
rect 3933 9131 4007 9145
rect 3727 9123 3761 9127
rect 3929 9115 4007 9131
rect 4073 9139 4147 9145
rect 4073 9134 4157 9139
rect 4073 9115 4147 9134
rect 3929 9111 3981 9115
rect 4181 9113 4287 9145
rect 4336 9135 4352 9139
rect 4371 9135 4405 9145
rect 4321 9111 4437 9135
rect 4458 9134 4479 9139
rect 4533 9134 4585 9139
rect 4591 9117 4593 9145
rect 4659 9117 4706 9145
rect 5107 9141 5449 9145
rect 5157 9134 5175 9137
rect 5239 9134 5266 9137
rect 5407 9134 5454 9137
rect 5491 9134 5543 9137
rect 3929 9084 3947 9097
rect 4321 9084 4437 9101
rect 3698 9080 5110 9084
rect 3929 9077 3947 9080
rect 4321 9077 4437 9080
rect 3670 9052 5082 9056
rect 13472 8986 13676 8988
rect 2044 8832 2310 8836
rect 2360 8832 3444 8836
rect 2044 8804 2310 8808
rect 2318 8806 2354 8816
rect 2360 8806 3416 8808
rect 2318 8804 3416 8806
rect 2280 8765 2283 8777
rect 2318 8772 2375 8804
rect 3386 8788 3416 8790
rect 3420 8788 3450 8824
rect 3574 8818 3576 8821
rect 3540 8784 3542 8788
rect 3574 8787 3623 8818
rect 2101 8743 2199 8763
rect 2249 8743 2283 8765
rect 2341 8743 2375 8772
rect 2407 8743 2486 8771
rect 2490 8767 2492 8781
rect 2793 8767 2796 8781
rect 2490 8763 2562 8767
rect 2584 8763 2670 8767
rect 2490 8749 2681 8763
rect 2683 8749 2796 8767
rect 2930 8761 2972 8767
rect 2920 8759 2972 8761
rect 2823 8749 2890 8759
rect 2919 8749 2972 8759
rect 2262 8739 2277 8743
rect 2066 8725 2096 8739
rect 2251 8735 2277 8739
rect 2101 8725 2199 8729
rect 2066 8713 2199 8725
rect 2067 8711 2199 8713
rect 2235 8713 2277 8735
rect 2235 8711 2279 8713
rect 2072 8709 2199 8711
rect 2072 8695 2174 8709
rect 2209 8701 2225 8711
rect 2235 8705 2273 8711
rect 2263 8701 2267 8705
rect 2219 8699 2225 8701
rect 2111 8691 2141 8695
rect 2072 8661 2084 8691
rect 2106 8684 2141 8691
rect 2096 8654 2141 8684
rect 2096 8644 2108 8654
rect 2120 8647 2140 8654
rect 2120 8644 2148 8647
rect 2096 8632 2148 8644
rect 2017 8629 2148 8632
rect 2054 8535 2066 8601
rect 2120 8589 2140 8629
rect 2154 8572 2174 8695
rect 2211 8673 2237 8699
rect 2195 8572 2200 8651
rect 2150 8556 2200 8572
rect 2195 8555 2200 8556
rect 2211 8647 2225 8673
rect 2269 8651 2273 8705
rect 2303 8669 2307 8743
rect 2354 8693 2368 8743
rect 2490 8739 2492 8749
rect 2520 8743 2596 8749
rect 2617 8743 2681 8749
rect 2682 8739 2683 8749
rect 2441 8713 2486 8737
rect 2532 8713 2534 8739
rect 2554 8713 2596 8729
rect 2646 8727 2647 8729
rect 2613 8713 2647 8727
rect 2724 8713 2725 8739
rect 2793 8713 2796 8749
rect 3019 8743 3131 8771
rect 3171 8749 3186 8767
rect 3192 8761 3258 8767
rect 3276 8765 3306 8767
rect 3261 8761 3306 8765
rect 3312 8761 3356 8767
rect 3192 8749 3356 8761
rect 3512 8750 3589 8784
rect 3555 8749 3589 8750
rect 3192 8743 3352 8749
rect 2441 8709 2647 8713
rect 2388 8693 2402 8709
rect 2478 8705 2647 8709
rect 2478 8701 2635 8705
rect 2478 8698 2507 8701
rect 2211 8566 2247 8647
rect 2326 8646 2454 8693
rect 2478 8647 2492 8698
rect 2554 8667 2635 8701
rect 2562 8657 2604 8667
rect 2373 8641 2454 8646
rect 2475 8641 2528 8647
rect 2373 8629 2448 8641
rect 2478 8629 2495 8641
rect 2562 8629 2640 8630
rect 2373 8612 2394 8629
rect 2211 8560 2225 8566
rect 2229 8560 2234 8566
rect 2211 8545 2240 8560
rect 2267 8545 2269 8583
rect 2263 8535 2269 8545
rect 2301 8535 2303 8549
rect 2475 8547 2494 8607
rect 2509 8555 2528 8613
rect 2646 8565 2647 8701
rect 2670 8698 2698 8713
rect 2670 8644 2683 8698
rect 2756 8675 2811 8713
rect 2819 8675 2821 8701
rect 2867 8690 2919 8705
rect 2793 8667 2811 8675
rect 2867 8667 2884 8690
rect 2787 8644 2884 8667
rect 2670 8629 2698 8644
rect 2778 8641 2884 8644
rect 2778 8633 2811 8641
rect 2680 8615 2681 8629
rect 2670 8599 2683 8615
rect 2670 8585 2718 8599
rect 2724 8585 2725 8629
rect 2753 8607 2840 8633
rect 2681 8581 2718 8585
rect 2681 8573 2726 8581
rect 2752 8573 2806 8599
rect 2712 8565 2726 8573
rect 2407 8535 2436 8547
rect 2441 8535 2475 8547
rect 2509 8535 2530 8555
rect 2647 8539 2726 8565
rect 2752 8539 2772 8565
rect 2712 8535 2726 8539
rect 2759 8535 2772 8539
rect 2793 8535 2806 8539
rect 2807 8535 2808 8607
rect 2890 8592 2919 8690
rect 3019 8675 3022 8743
rect 3035 8739 3050 8743
rect 3035 8737 3061 8739
rect 3117 8737 3138 8739
rect 3035 8713 3138 8737
rect 3192 8713 3198 8743
rect 3216 8717 3222 8739
rect 3226 8713 3318 8727
rect 3326 8713 3352 8743
rect 3053 8709 3131 8713
rect 3053 8675 3056 8709
rect 3087 8665 3088 8709
rect 3171 8698 3198 8713
rect 3221 8701 3368 8713
rect 3186 8669 3198 8698
rect 3226 8669 3232 8701
rect 3243 8698 3368 8701
rect 3186 8666 3192 8669
rect 3258 8667 3352 8698
rect 2920 8650 3053 8657
rect 3087 8650 3108 8665
rect 3180 8657 3232 8666
rect 2920 8641 3108 8650
rect 3011 8634 3016 8641
rect 2938 8623 3019 8634
rect 3046 8623 3108 8641
rect 3167 8635 3232 8657
rect 3258 8651 3292 8667
rect 3306 8651 3312 8667
rect 2920 8620 3108 8623
rect 2920 8607 3053 8620
rect 2875 8586 2919 8592
rect 2938 8587 3019 8607
rect 2867 8579 2970 8586
rect 2975 8579 3019 8587
rect 3125 8579 3141 8589
rect 2867 8577 3163 8579
rect 2893 8574 3163 8577
rect 3167 8574 3175 8623
rect 3186 8622 3192 8635
rect 3214 8622 3232 8632
rect 3271 8622 3292 8651
rect 3326 8633 3352 8667
rect 3305 8622 3326 8633
rect 3182 8596 3326 8622
rect 3356 8599 3368 8698
rect 3339 8596 3368 8599
rect 3555 8712 3578 8749
rect 3555 8596 3589 8712
rect 3182 8575 3368 8596
rect 3201 8574 3209 8575
rect 1991 8531 2066 8535
rect 2073 8531 2362 8535
rect 1991 8521 2362 8531
rect 1991 8497 2066 8521
rect 2073 8497 2362 8521
rect 2407 8523 2598 8535
rect 2621 8523 2731 8535
rect 2759 8531 2878 8535
rect 2407 8515 2731 8523
rect 1991 8493 2362 8497
rect 2412 8493 2731 8515
rect 2761 8515 2878 8531
rect 2893 8515 3214 8574
rect 2761 8513 3214 8515
rect 3222 8557 3368 8575
rect 3512 8593 3589 8596
rect 3222 8535 3292 8557
rect 3305 8549 3368 8557
rect 3305 8535 3326 8549
rect 3339 8535 3368 8549
rect 3373 8535 3394 8565
rect 3512 8562 3541 8593
rect 3555 8573 3589 8593
rect 3544 8562 3589 8573
rect 3595 8535 3623 8595
rect 3862 8542 3904 8552
rect 3864 8538 3904 8542
rect 3222 8525 3652 8535
rect 3222 8513 3264 8525
rect 2737 8493 2752 8509
rect 2761 8493 3180 8513
rect 3192 8511 3219 8513
rect 3190 8493 3219 8511
rect 3271 8512 3652 8525
rect 3834 8514 3876 8524
rect 3271 8493 3650 8512
rect 3836 8510 3876 8514
rect 1991 8488 3650 8493
rect 1991 8477 3454 8488
rect 2111 8467 2138 8477
rect 2151 8467 2183 8477
rect 2195 8467 2200 8477
rect 2229 8467 2234 8477
rect 2059 8463 2111 8467
rect 2141 8463 2234 8467
rect 2059 8453 2195 8463
rect 2059 8429 2137 8453
rect 2141 8452 2195 8453
rect 2151 8429 2195 8452
rect 2229 8455 2234 8463
rect 2059 8417 2201 8429
rect 2059 8391 2161 8417
rect 2041 8387 2161 8391
rect 1998 8383 2161 8387
rect 1998 8369 2163 8383
rect 2111 8357 2127 8369
rect 2135 8357 2163 8369
rect 2135 8353 2161 8357
rect 2177 8353 2201 8417
rect 2229 8383 2235 8455
rect 2267 8405 2269 8477
rect 2271 8383 2277 8445
rect 2301 8387 2303 8477
rect 2447 8467 2480 8477
rect 2347 8465 2477 8467
rect 2347 8452 2362 8465
rect 2367 8455 2477 8465
rect 2383 8453 2477 8455
rect 2309 8387 2315 8407
rect 2345 8398 2381 8445
rect 2395 8421 2477 8453
rect 2481 8431 2509 8477
rect 2737 8467 2752 8477
rect 2771 8467 2806 8475
rect 2511 8455 2530 8467
rect 2689 8457 2806 8467
rect 2671 8455 2806 8457
rect 2840 8467 2938 8477
rect 2961 8467 3011 8477
rect 2840 8455 3011 8467
rect 2511 8440 2641 8455
rect 2511 8429 2621 8440
rect 2395 8405 2449 8421
rect 2515 8409 2545 8429
rect 2395 8401 2425 8405
rect 2491 8401 2545 8409
rect 2549 8423 2621 8429
rect 2635 8423 2641 8440
rect 2645 8452 2786 8455
rect 2863 8452 2879 8455
rect 2645 8423 2717 8452
rect 2549 8401 2689 8423
rect 2731 8401 2761 8452
rect 2771 8401 2786 8452
rect 2878 8415 2879 8452
rect 2888 8431 3011 8455
rect 2909 8415 3011 8431
rect 3035 8476 3112 8477
rect 3035 8464 3114 8476
rect 2919 8401 2949 8415
rect 2395 8398 2964 8401
rect 2211 8353 2235 8383
rect 2301 8357 2341 8387
rect 2345 8383 2964 8398
rect 3001 8387 3006 8415
rect 3035 8391 3040 8464
rect 3041 8455 3107 8464
rect 3180 8455 3182 8477
rect 3271 8467 3292 8477
rect 3305 8467 3345 8477
rect 3373 8475 3394 8477
rect 3265 8465 3326 8467
rect 3041 8415 3110 8455
rect 3165 8443 3224 8455
rect 3249 8443 3326 8465
rect 3165 8440 3306 8443
rect 13472 8442 13477 8476
rect 13472 8441 13511 8442
rect 3180 8431 3306 8440
rect 3180 8415 3219 8431
rect 3249 8415 3306 8431
rect 3041 8393 3046 8415
rect 3108 8393 3110 8415
rect 3055 8391 3089 8393
rect 3149 8387 3258 8415
rect 3276 8393 3306 8415
rect 3339 8393 3360 8421
rect 2407 8357 2447 8383
rect 2450 8357 2467 8383
rect 2491 8379 2522 8383
rect 2549 8379 2655 8383
rect 2491 8357 2521 8379
rect 2545 8363 2655 8379
rect 2689 8369 2723 8383
rect 2771 8363 2786 8383
rect 2545 8357 2621 8363
rect 2919 8359 2949 8383
rect 2993 8359 3006 8387
rect 3276 8383 3291 8393
rect 2549 8355 2621 8357
rect 2893 8357 2959 8359
rect 3011 8357 3016 8383
rect 3138 8357 3140 8383
rect 3222 8381 3249 8383
rect 2893 8353 2925 8357
rect 2927 8353 2959 8357
rect 3148 8353 3182 8381
rect 3216 8353 3258 8381
rect 3315 8357 3360 8393
rect 3339 8353 3360 8357
rect 3373 8353 3394 8436
rect 3411 8391 3464 8414
rect 3404 8383 3464 8391
rect 3494 8411 3585 8414
rect 3494 8383 3604 8411
rect 3458 8358 3550 8360
rect 3458 8357 3505 8358
rect 2032 8335 2161 8353
rect 2267 8339 2341 8353
rect 2061 8331 2095 8335
rect 2263 8323 2341 8339
rect 2407 8347 2481 8353
rect 2407 8342 2491 8347
rect 2407 8323 2481 8342
rect 2263 8319 2315 8323
rect 2515 8321 2621 8353
rect 2670 8343 2686 8347
rect 2705 8343 2739 8353
rect 2655 8319 2771 8343
rect 2792 8342 2813 8347
rect 2867 8342 2919 8347
rect 2925 8325 2927 8353
rect 2993 8325 3040 8353
rect 3458 8349 3464 8357
rect 3494 8349 3505 8357
rect 3544 8346 3550 8358
rect 2263 8292 2281 8305
rect 2655 8292 2771 8309
rect 2032 8288 3780 8292
rect 2263 8285 2281 8288
rect 2655 8285 2771 8288
rect 8184 8272 11394 8306
rect 2004 8260 3752 8264
rect 1966 8168 2876 8190
rect 2692 8162 2804 8168
rect 1966 8140 2876 8162
rect 4506 8156 4652 8192
rect 7464 8156 7498 8212
rect 7643 8160 7851 8190
rect 7647 8156 7810 8160
rect 7846 8156 7847 8160
rect 7996 8156 8030 8212
rect 8088 8156 8122 8210
rect 9853 8204 9854 8258
rect 8267 8158 9014 8190
rect 9907 8183 9908 8204
rect 9919 8183 11295 8192
rect 2024 8076 2502 8084
rect 2692 8082 2804 8140
rect 2574 8080 2976 8082
rect 2574 8076 2944 8080
rect 1054 8042 1056 8052
rect 2052 8048 2502 8056
rect 2692 8054 2804 8076
rect 2574 8048 2948 8054
rect 1026 8014 1056 8024
rect 2692 7890 2804 8048
rect 2913 8019 2955 8031
rect 2879 7985 2985 7997
rect 2995 7933 2999 7959
rect 3079 7933 3107 7959
rect 3005 7921 3039 7933
rect 3133 7931 3149 7933
rect 3005 7899 3047 7921
rect 2703 7889 2804 7890
rect 3013 7887 3047 7899
rect 3049 7887 3057 7931
rect 3133 7887 3161 7931
rect 3173 7917 3185 7933
rect 3173 7899 3215 7917
rect 3185 7891 3215 7899
rect 3223 7913 3257 7917
rect 3269 7913 3299 7917
rect 3223 7899 3299 7913
rect 3223 7895 3257 7899
rect 3269 7891 3299 7899
rect 2939 7787 2955 7883
rect 2965 7880 2969 7881
rect 2973 7880 2989 7883
rect 3133 7881 3149 7887
rect 3185 7881 3205 7891
rect 3049 7880 3077 7881
rect 3133 7880 3163 7881
rect 3217 7880 3247 7891
rect 3269 7881 3289 7891
rect 2958 7849 3013 7880
rect 3042 7849 3117 7880
rect 3126 7849 3346 7880
rect 2958 7833 3346 7849
rect 2965 7787 2969 7833
rect 2973 7787 2989 7833
rect 2999 7819 3077 7833
rect 3089 7823 3346 7833
rect 3089 7819 3433 7823
rect 2999 7815 3433 7819
rect 3650 7817 3828 8138
rect 4506 8122 8980 8156
rect 4506 7832 4652 8122
rect 7430 7933 7442 7999
rect 4506 7831 4645 7832
rect 4506 7817 4532 7831
rect 2999 7807 3499 7815
rect 7464 7810 7498 8122
rect 7571 8054 7600 8080
rect 7571 8042 7647 8054
rect 7847 8042 7959 8054
rect 7996 8042 8030 8122
rect 7571 8039 7959 8042
rect 7571 8033 7944 8039
rect 7566 8008 7944 8033
rect 7962 8008 8030 8042
rect 7516 7933 7550 7999
rect 7566 7996 7647 8008
rect 7847 7996 7944 8008
rect 7566 7970 7600 7996
rect 7566 7962 7588 7970
rect 7597 7962 7600 7970
rect 7566 7936 7600 7962
rect 7894 7937 7928 7996
rect 7847 7936 7928 7937
rect 7566 7924 7647 7936
rect 7847 7924 7944 7936
rect 7996 7924 8030 8008
rect 8088 8042 8122 8122
rect 8190 8099 8224 8101
rect 8946 8074 8980 8122
rect 8283 8042 8980 8074
rect 9820 8149 9831 8160
rect 9843 8149 9854 8160
rect 9903 8158 11311 8183
rect 11352 8160 11361 8258
rect 9907 8152 9992 8158
rect 11203 8152 11307 8158
rect 9907 8149 9956 8152
rect 11203 8150 11284 8152
rect 11203 8149 11298 8150
rect 11352 8149 11363 8160
rect 11375 8149 11386 8160
rect 9820 8083 9854 8149
rect 9906 8146 9972 8149
rect 11203 8146 11300 8149
rect 9879 8124 9964 8146
rect 11203 8133 11298 8146
rect 11352 8145 11386 8149
rect 11242 8124 11298 8133
rect 11348 8133 11394 8145
rect 9922 8108 9956 8124
rect 11250 8108 11284 8124
rect 9820 8072 9831 8083
rect 9843 8072 9854 8083
rect 9879 8086 9964 8108
rect 11242 8086 11298 8108
rect 11348 8099 11386 8133
rect 11348 8087 11394 8099
rect 8088 8040 8980 8042
rect 8088 8008 8785 8040
rect 8797 8028 8925 8030
rect 8088 7960 8122 8008
rect 8844 7983 8878 7994
rect 8946 7960 8980 8040
rect 9879 8006 9890 8086
rect 9906 8083 9972 8086
rect 11234 8083 11300 8086
rect 11352 8083 11386 8087
rect 9907 8080 9922 8083
rect 11242 8082 11298 8083
rect 9907 8074 9992 8080
rect 11214 8074 11307 8080
rect 9903 8049 11311 8074
rect 11352 8072 11363 8083
rect 11375 8072 11386 8083
rect 9907 8034 9918 8049
rect 9919 8040 11295 8049
rect 9907 8028 9908 8034
rect 11352 8028 11361 8072
rect 8088 7926 11394 7960
rect 7566 7899 7944 7924
rect 7571 7893 7944 7899
rect 7962 7910 8030 7924
rect 8054 7910 8801 7924
rect 7571 7890 7959 7893
rect 7962 7892 8801 7910
rect 7962 7890 8797 7892
rect 7571 7878 7647 7890
rect 7847 7878 7959 7890
rect 7968 7886 8797 7890
rect 8946 7886 8980 7926
rect 7968 7884 9016 7886
rect 7996 7882 8030 7884
rect 8052 7882 9016 7884
rect 7571 7852 7600 7878
rect 7996 7856 9016 7882
rect 7996 7810 8030 7856
rect 8044 7810 8064 7828
rect 8070 7810 9016 7856
rect 2999 7799 3285 7807
rect 3302 7806 3499 7807
rect 3302 7799 3315 7806
rect 2999 7787 3077 7799
rect 3107 7787 3285 7799
rect 2826 7750 2868 7768
rect 2887 7750 3325 7787
rect 3336 7772 3399 7789
rect 3456 7772 3499 7781
rect 4638 7776 9016 7810
rect 3336 7765 3349 7772
rect 2716 7700 2736 7726
rect 2750 7700 2770 7734
rect 2826 7697 3325 7750
rect 7464 7706 7498 7776
rect 7566 7748 7600 7776
rect 7894 7748 7928 7776
rect 7996 7706 8030 7776
rect 8044 7706 8064 7776
rect 8070 7740 9016 7776
rect 8070 7706 8604 7740
rect 2868 7695 2973 7696
rect 2995 7685 3215 7697
rect 3268 7685 3299 7697
rect 2995 7667 3055 7685
rect 2839 7613 2842 7667
rect 2913 7631 2965 7667
rect 2969 7635 3055 7667
rect 3057 7677 3129 7685
rect 3057 7667 3107 7677
rect 3115 7667 3123 7677
rect 3057 7635 3133 7667
rect 3149 7660 3157 7685
rect 3163 7660 3215 7685
rect 3138 7649 3230 7660
rect 3269 7649 3299 7685
rect 5262 7672 8604 7706
rect 3138 7642 3299 7649
rect 3154 7640 3299 7642
rect 3157 7635 3299 7640
rect 2969 7631 3049 7635
rect 3077 7632 3133 7635
rect 3159 7632 3299 7635
rect 3077 7631 3299 7632
rect 2919 7613 2969 7631
rect 2893 7552 2896 7613
rect 2939 7605 2969 7613
rect 2939 7601 2965 7605
rect 2973 7601 2989 7631
rect 3027 7613 3077 7631
rect 3034 7605 3077 7613
rect 2950 7598 2965 7601
rect 3034 7598 3049 7605
rect 3081 7601 3089 7631
rect 3110 7614 3258 7631
rect 3123 7613 3257 7614
rect 3118 7601 3257 7613
rect 3269 7605 3289 7631
rect 3118 7598 3133 7601
rect 3144 7595 3159 7601
rect 3144 7590 3178 7595
rect 3215 7590 3262 7595
rect 3023 7567 3201 7579
rect 2876 7536 2972 7538
rect 3023 7533 3083 7545
rect 3117 7533 3167 7545
rect 2848 7508 2944 7510
rect 2460 7396 2502 7414
rect 2574 7396 3662 7414
rect 2864 7392 3662 7396
rect 2864 7388 3416 7392
rect 2432 7368 2502 7386
rect 2574 7368 3662 7386
rect 2836 7364 3662 7368
rect 2836 7360 3444 7364
rect 2022 7290 2293 7294
rect 2358 7290 3434 7294
rect 3350 7266 3376 7272
rect 1994 7262 2293 7266
rect 2306 7258 2346 7266
rect 2358 7262 3406 7266
rect 2268 7223 2273 7235
rect 2306 7224 2365 7258
rect 1227 7219 1261 7223
rect 786 7038 844 7206
rect 1198 7201 1301 7219
rect 1319 7201 1353 7223
rect 1367 7201 1410 7219
rect 2091 7201 2189 7221
rect 2239 7201 2273 7223
rect 2331 7201 2365 7224
rect 2397 7201 2476 7229
rect 2480 7225 2482 7239
rect 2783 7225 2786 7239
rect 3350 7235 3376 7262
rect 3384 7235 3410 7238
rect 3460 7235 3490 7238
rect 3494 7235 3524 7269
rect 3564 7245 3571 7269
rect 2480 7221 2552 7225
rect 2574 7221 2660 7225
rect 2480 7207 2671 7221
rect 2673 7207 2786 7225
rect 2920 7219 2962 7225
rect 2910 7217 2962 7219
rect 2813 7207 2880 7217
rect 2909 7207 2962 7217
rect 2252 7197 2267 7201
rect 2056 7196 2086 7197
rect 1164 7167 1301 7185
rect 1221 7163 1255 7167
rect 1313 7163 1347 7185
rect 1367 7151 1376 7185
rect 1386 7170 1469 7196
rect 1534 7170 2213 7196
rect 2241 7193 2267 7197
rect 2225 7171 2267 7193
rect 2057 7169 2189 7170
rect 2225 7169 2269 7171
rect 2062 7168 2189 7169
rect 2199 7168 2215 7169
rect 1241 7143 1271 7147
rect 1233 7121 1271 7143
rect 1301 7121 1351 7135
rect 1233 7117 1267 7121
rect 1199 7083 1227 7109
rect 1277 7101 1351 7121
rect 1401 7117 1410 7167
rect 1414 7142 1469 7168
rect 1534 7157 2215 7168
rect 2225 7157 2263 7169
rect 1534 7151 2263 7157
rect 1444 7103 1477 7137
rect 1482 7104 1522 7146
rect 1534 7142 2227 7151
rect 2086 7137 2131 7142
rect 2144 7137 2164 7142
rect 2201 7137 2227 7142
rect 2259 7137 2263 7151
rect 2293 7137 2297 7201
rect 2344 7151 2358 7201
rect 2480 7197 2482 7207
rect 2510 7201 2586 7207
rect 2607 7201 2671 7207
rect 2672 7197 2673 7207
rect 2431 7171 2476 7195
rect 2522 7171 2524 7197
rect 2544 7171 2586 7187
rect 2636 7185 2637 7187
rect 2603 7171 2637 7185
rect 2714 7171 2715 7197
rect 2783 7171 2786 7207
rect 3009 7201 3121 7229
rect 3161 7207 3176 7225
rect 3182 7219 3248 7225
rect 3266 7223 3296 7225
rect 3251 7219 3296 7223
rect 3302 7219 3346 7225
rect 3182 7207 3346 7219
rect 3460 7207 3537 7235
rect 3182 7201 3342 7207
rect 3460 7201 3495 7207
rect 2431 7167 2637 7171
rect 2378 7151 2392 7167
rect 2468 7159 2637 7167
rect 2468 7156 2497 7159
rect 1535 7103 1560 7137
rect 2062 7127 2144 7137
rect 1738 7123 1750 7127
rect 1761 7123 1819 7127
rect 1576 7109 1628 7121
rect 1658 7117 1702 7121
rect 1573 7103 1652 7109
rect 1241 7083 1267 7093
rect 1233 7067 1267 7083
rect 1277 7075 1335 7101
rect 1414 7090 1475 7099
rect 1573 7090 1628 7103
rect 1658 7090 1713 7117
rect 1738 7101 1819 7123
rect 1844 7115 1966 7127
rect 1989 7119 2144 7127
rect 2187 7131 2227 7137
rect 1989 7115 2065 7119
rect 1844 7103 2065 7115
rect 1233 7051 1271 7067
rect 1277 7051 1307 7075
rect 1414 7072 1734 7090
rect 1738 7087 1834 7101
rect 1844 7090 1966 7103
rect 1989 7092 2065 7103
rect 2086 7092 2138 7119
rect 2187 7113 2215 7131
rect 2271 7113 2297 7137
rect 2201 7103 2215 7113
rect 2278 7103 2297 7109
rect 2316 7104 2444 7151
rect 2468 7127 2482 7156
rect 2544 7151 2637 7159
rect 2468 7105 2522 7127
rect 2544 7125 2625 7151
rect 2636 7137 2637 7151
rect 2660 7156 2688 7171
rect 2739 7167 2740 7171
rect 2660 7137 2673 7156
rect 2639 7127 2673 7137
rect 2705 7133 2740 7137
rect 2746 7133 2801 7171
rect 2809 7167 2865 7171
rect 2910 7167 2944 7171
rect 2857 7148 2909 7163
rect 2783 7127 2801 7133
rect 2639 7125 2714 7127
rect 2738 7125 2801 7127
rect 2804 7137 2838 7141
rect 2857 7137 2874 7148
rect 2804 7133 2874 7137
rect 2552 7115 2598 7125
rect 2565 7113 2598 7115
rect 2639 7113 2802 7125
rect 2568 7105 2598 7113
rect 1989 7090 2138 7092
rect 2144 7090 2164 7103
rect 2178 7090 2190 7103
rect 2201 7090 2224 7103
rect 2263 7090 2278 7103
rect 2297 7099 2312 7103
rect 2283 7090 2312 7099
rect 2337 7090 2352 7104
rect 2363 7099 2444 7104
rect 2465 7099 2522 7105
rect 2552 7103 2598 7105
rect 2654 7103 2802 7113
rect 2568 7102 2598 7103
rect 2363 7090 2522 7099
rect 1844 7087 2522 7090
rect 2553 7087 2613 7102
rect 2636 7087 2637 7103
rect 2654 7091 2714 7103
rect 2738 7099 2802 7103
rect 2804 7099 2838 7133
rect 2857 7099 2874 7133
rect 2880 7099 2909 7148
rect 3009 7137 3012 7201
rect 3025 7197 3040 7201
rect 3025 7195 3051 7197
rect 3107 7195 3128 7197
rect 3025 7171 3128 7195
rect 3182 7171 3188 7201
rect 3206 7175 3212 7197
rect 3316 7196 3342 7201
rect 3273 7185 3406 7196
rect 3216 7171 3406 7185
rect 3043 7167 3122 7171
rect 3043 7137 3046 7167
rect 3077 7161 3122 7167
rect 3077 7137 3078 7161
rect 3161 7156 3188 7171
rect 3211 7170 3406 7171
rect 3527 7170 3537 7207
rect 3211 7168 3358 7170
rect 3211 7159 3434 7168
rect 3176 7137 3188 7156
rect 3216 7137 3222 7159
rect 3227 7151 3434 7159
rect 3248 7142 3434 7151
rect 3248 7137 3342 7142
rect 3346 7141 3358 7142
rect 2910 7133 2944 7137
rect 3077 7127 3122 7137
rect 3077 7123 3078 7127
rect 3077 7115 3098 7123
rect 2910 7099 2956 7115
rect 3025 7108 3043 7115
rect 3077 7108 3115 7115
rect 2738 7091 2801 7099
rect 2654 7087 2802 7091
rect 1813 7073 1834 7087
rect 1415 7071 1435 7072
rect 1233 7049 1307 7051
rect 1267 7033 1307 7049
rect 1389 7062 1447 7071
rect 1573 7062 1583 7072
rect 1607 7069 1652 7072
rect 1607 7067 1617 7069
rect 1628 7067 1649 7069
rect 1607 7062 1659 7067
rect 1686 7066 1719 7072
rect 1389 7048 1734 7062
rect 1792 7055 1801 7073
rect 1804 7058 1844 7073
rect 1813 7055 1844 7058
rect 1386 7044 1734 7048
rect 1277 7022 1307 7033
rect 1271 7017 1307 7022
rect 807 6983 938 7011
rect 971 6995 1193 7007
rect 1267 6999 1307 7017
rect 1031 6983 1193 6995
rect 1271 6992 1307 6999
rect 1346 6994 1347 7037
rect 1401 7031 1435 7044
rect 1573 7031 1583 7044
rect 1607 7031 1617 7044
rect 1493 7019 1617 7031
rect 1628 7041 1685 7044
rect 1271 6983 1274 6992
rect 1336 6985 1347 6994
rect 1363 6993 1389 7017
rect 1447 6993 1473 7017
rect 1492 7000 1620 7019
rect 1628 7017 1658 7041
rect 1779 7031 1844 7055
rect 1628 7007 1685 7017
rect 1628 7005 1658 7007
rect 1628 7000 1665 7005
rect 1285 6983 1347 6985
rect 1492 6985 1665 7000
rect 1704 6995 1770 7021
rect 1792 7011 1801 7031
rect 1813 7017 1844 7031
rect 1847 7017 1868 7087
rect 1934 7083 2479 7087
rect 2522 7083 2541 7087
rect 2568 7083 2594 7087
rect 1884 7069 1915 7081
rect 1934 7076 2594 7083
rect 2630 7076 2640 7087
rect 2670 7076 2671 7087
rect 2705 7076 2810 7087
rect 1934 7074 2826 7076
rect 2831 7074 2909 7099
rect 2939 7081 2960 7099
rect 2910 7074 2960 7081
rect 3001 7092 3006 7108
rect 3025 7103 3115 7108
rect 3025 7099 3098 7103
rect 3009 7092 3025 7099
rect 3036 7092 3098 7099
rect 3157 7093 3160 7115
rect 3176 7093 3182 7137
rect 3191 7113 3225 7137
rect 3248 7125 3339 7137
rect 3248 7109 3316 7125
rect 3261 7103 3316 7109
rect 3001 7081 3098 7092
rect 3126 7081 3157 7093
rect 3160 7083 3191 7093
rect 3222 7083 3252 7099
rect 3261 7083 3282 7103
rect 3346 7099 3376 7141
rect 3454 7109 3470 7141
rect 3526 7120 3537 7170
rect 4506 7176 4668 7648
rect 6931 7604 6932 7658
rect 6957 7604 7120 7626
rect 7560 7622 7934 7626
rect 8010 7604 8030 7672
rect 6985 7598 6986 7604
rect 6985 7592 7148 7598
rect 7464 7592 8030 7604
rect 8044 7592 8064 7672
rect 8070 7592 8604 7672
rect 9402 7626 9658 7630
rect 9430 7598 9630 7602
rect 6985 7583 8604 7592
rect 6898 7549 6909 7560
rect 6921 7549 6932 7560
rect 6981 7558 8604 7583
rect 6985 7552 7070 7558
rect 6985 7549 7034 7552
rect 6898 7483 6932 7549
rect 6984 7546 7050 7549
rect 6957 7524 7042 7546
rect 7000 7508 7034 7524
rect 6898 7472 6909 7483
rect 6921 7472 6932 7483
rect 6957 7486 7042 7508
rect 6957 7424 6968 7486
rect 6984 7483 7050 7486
rect 6985 7480 7000 7483
rect 6985 7474 7070 7480
rect 8070 7474 8604 7558
rect 6981 7449 8604 7474
rect 6985 7440 8604 7449
rect 6985 7434 7206 7440
rect 7266 7434 8604 7440
rect 9676 7436 9769 7439
rect 9676 7435 9808 7436
rect 6985 7428 6986 7434
rect 8070 7424 8604 7434
rect 9660 7432 9808 7435
rect 9944 7433 9964 7436
rect 6957 7406 7206 7424
rect 7266 7406 8604 7424
rect 8070 7360 8604 7406
rect 5262 7326 8604 7360
rect 8070 7290 8604 7326
rect 9262 7420 9798 7422
rect 9944 7420 9978 7433
rect 9262 7282 10008 7420
rect 9262 7266 9462 7282
rect 4506 7152 4686 7176
rect 9020 7174 9048 7176
rect 4506 7148 4668 7152
rect 4506 7124 4714 7148
rect 3503 7109 3514 7110
rect 3409 7103 3514 7109
rect 3314 7091 3344 7099
rect 3346 7091 3358 7099
rect 3295 7083 3358 7091
rect 3160 7081 3358 7083
rect 3001 7078 3115 7081
rect 3001 7074 3056 7078
rect 3077 7074 3115 7078
rect 3128 7074 3155 7081
rect 3157 7074 3160 7081
rect 3176 7080 3182 7081
rect 3187 7080 3358 7081
rect 3172 7074 3358 7080
rect 1934 7073 3358 7074
rect 3398 7078 3418 7099
rect 3454 7078 3470 7103
rect 3503 7099 3514 7103
rect 3526 7109 3545 7120
rect 3503 7095 3512 7099
rect 3526 7095 3537 7109
rect 3503 7078 3537 7095
rect 3398 7073 3537 7078
rect 3551 7073 3566 7087
rect 1934 7072 3391 7073
rect 3403 7072 3574 7073
rect 1949 7069 2190 7072
rect 1966 7062 2004 7069
rect 2007 7062 2190 7069
rect 2201 7062 2224 7072
rect 2278 7069 2297 7072
rect 2337 7062 2354 7072
rect 2371 7071 2397 7072
rect 2405 7071 2568 7072
rect 2371 7065 2569 7071
rect 2598 7069 2654 7072
rect 2670 7070 2671 7072
rect 2699 7070 2852 7072
rect 2391 7062 2569 7065
rect 1934 7058 2569 7062
rect 1934 7055 2518 7058
rect 2522 7055 2569 7058
rect 1934 7053 2569 7055
rect 1922 7051 2569 7053
rect 1918 7048 2569 7051
rect 2594 7048 2654 7069
rect 2665 7065 2852 7070
rect 2665 7061 2842 7065
rect 2665 7058 2836 7061
rect 2665 7051 2793 7058
rect 2665 7048 2796 7051
rect 2797 7048 2827 7058
rect 2865 7049 2909 7072
rect 2910 7065 2956 7072
rect 3001 7061 3056 7072
rect 3077 7069 3115 7072
rect 3128 7065 3155 7072
rect 1918 7047 2827 7048
rect 1922 7046 2827 7047
rect 2880 7046 2918 7049
rect 2965 7047 3056 7061
rect 3098 7047 3125 7063
rect 3157 7059 3160 7072
rect 3172 7061 3391 7072
rect 2965 7046 3077 7047
rect 3081 7046 3125 7047
rect 3172 7057 3344 7061
rect 3346 7058 3388 7061
rect 3439 7058 3574 7072
rect 3626 7059 3654 7123
rect 4028 7101 4072 7123
rect 3660 7059 3688 7089
rect 3346 7057 3384 7058
rect 3172 7054 3404 7057
rect 3172 7053 3428 7054
rect 3172 7051 3438 7053
rect 3454 7051 3540 7058
rect 3172 7050 3444 7051
rect 3449 7050 3540 7051
rect 3172 7046 3540 7050
rect 1922 7044 3540 7046
rect 1815 7011 1849 7017
rect 1789 7007 1849 7011
rect 1872 7007 1874 7021
rect 1922 7017 2190 7044
rect 2201 7017 2224 7044
rect 2253 7041 2272 7044
rect 2278 7041 2305 7044
rect 2253 7017 2278 7041
rect 2305 7017 2312 7041
rect 1918 7015 2178 7017
rect 1918 7014 2175 7015
rect 1918 7013 2164 7014
rect 1966 7009 2135 7013
rect 1966 7007 2125 7009
rect 1741 6993 1757 6995
rect 1789 6989 1860 7007
rect 1872 7003 1944 7007
rect 1966 7003 2175 7007
rect 2183 7004 2216 7017
rect 2278 7007 2305 7017
rect 2352 7013 2354 7044
rect 2403 7043 2654 7044
rect 2403 7038 2603 7043
rect 2630 7038 2654 7043
rect 2665 7038 2796 7044
rect 2403 7031 2796 7038
rect 2797 7031 2827 7044
rect 2880 7037 2960 7044
rect 2965 7037 3077 7044
rect 2356 7017 2382 7021
rect 2424 7017 2793 7031
rect 2796 7028 2827 7031
rect 2830 7028 2852 7031
rect 2880 7028 3077 7037
rect 3081 7032 3125 7044
rect 3172 7033 3444 7044
rect 3182 7032 3444 7033
rect 3081 7028 3444 7032
rect 2796 7018 3444 7028
rect 2796 7017 2827 7018
rect 2356 7013 2401 7017
rect 2352 7007 2401 7013
rect 2183 7003 2230 7004
rect 2238 7003 2253 7004
rect 1872 7000 2178 7003
rect 1872 6989 2063 7000
rect 2065 6989 2178 7000
rect 1492 6984 1685 6985
rect 1529 6983 1685 6984
rect 1789 6983 1847 6989
rect 841 6949 904 6977
rect 1112 6973 1133 6979
rect 1031 6960 1159 6973
rect 1211 6972 1241 6979
rect 1267 6972 1347 6983
rect 1166 6963 1347 6972
rect 1354 6963 1366 6983
rect 1388 6963 1400 6983
rect 1166 6960 1400 6963
rect 1031 6954 1400 6960
rect 1448 6954 1478 6979
rect 1529 6969 1577 6983
rect 1581 6969 1659 6983
rect 1529 6963 1659 6969
rect 1685 6963 1689 6983
rect 1736 6963 1750 6983
rect 1529 6954 1761 6963
rect 807 6851 827 6949
rect 841 6851 861 6949
rect 968 6938 986 6953
rect 1031 6952 1761 6954
rect 1779 6953 1784 6983
rect 1789 6953 1813 6983
rect 1872 6979 1874 6989
rect 1902 6983 1978 6989
rect 1953 6979 1978 6983
rect 1980 6979 2063 6989
rect 2064 6979 2131 6989
rect 1823 6953 1847 6977
rect 1914 6953 1916 6979
rect 1936 6963 1978 6969
rect 2006 6967 2056 6979
rect 2106 6970 2136 6979
rect 1995 6963 2056 6967
rect 1936 6955 2045 6963
rect 1936 6954 2063 6955
rect 2097 6954 2131 6955
rect 2175 6954 2178 6989
rect 2183 6989 2272 7003
rect 2312 7001 2401 7007
rect 2302 6999 2401 7001
rect 2301 6993 2401 6999
rect 2424 7004 2796 7017
rect 2797 7004 2827 7017
rect 2830 7011 2852 7018
rect 2880 7017 3444 7018
rect 2880 7013 3204 7017
rect 2424 7000 2842 7004
rect 2876 7000 3204 7013
rect 3212 7015 3444 7017
rect 3212 7000 3282 7015
rect 3295 7000 3444 7015
rect 2424 6997 3444 7000
rect 2424 6994 2499 6997
rect 2301 6989 2382 6993
rect 2183 6983 2216 6989
rect 2230 6973 2249 6989
rect 2253 6988 2257 6989
rect 2352 6979 2382 6989
rect 2417 6989 2499 6994
rect 2417 6983 2432 6989
rect 2440 6983 2499 6989
rect 2512 6989 3444 6997
rect 2512 6983 2598 6989
rect 2608 6983 2736 6989
rect 2745 6983 2886 6989
rect 2215 6958 2272 6973
rect 2352 6963 2373 6979
rect 2397 6977 2469 6983
rect 2512 6979 2553 6983
rect 2499 6977 2553 6979
rect 2397 6963 2553 6977
rect 2230 6954 2249 6958
rect 2352 6954 2553 6963
rect 1934 6953 2553 6954
rect 2568 6979 2598 6983
rect 2603 6979 2646 6983
rect 2568 6975 2646 6979
rect 2568 6957 2658 6975
rect 2702 6973 2736 6983
rect 2568 6953 2653 6957
rect 2674 6955 2700 6967
rect 2708 6955 2736 6973
rect 2674 6953 2708 6955
rect 2721 6953 2736 6955
rect 2749 6981 2886 6983
rect 2925 6983 3444 6989
rect 3449 7001 3540 7044
rect 3449 6985 3498 7001
rect 2925 6981 3296 6983
rect 2749 6953 2909 6981
rect 1031 6949 1159 6952
rect 1050 6938 1070 6949
rect 1143 6939 1163 6949
rect 968 6923 971 6938
rect 960 6920 1010 6923
rect 1050 6920 1055 6938
rect 1091 6920 1094 6939
rect 1125 6932 1128 6939
rect 1153 6932 1163 6939
rect 1183 6932 1366 6952
rect 1110 6926 1366 6932
rect 1381 6938 1406 6952
rect 1449 6951 1478 6952
rect 1493 6939 1520 6951
rect 1529 6950 1761 6952
rect 1529 6949 1581 6950
rect 1529 6939 1577 6949
rect 1591 6941 1761 6950
rect 1774 6949 1847 6953
rect 1860 6951 2499 6953
rect 2520 6951 2580 6953
rect 2603 6951 2909 6953
rect 2925 6971 3204 6981
rect 3212 6971 3239 6981
rect 3266 6971 3294 6981
rect 3305 6973 3444 6983
rect 3305 6971 3407 6973
rect 2925 6951 3222 6971
rect 3266 6951 3296 6971
rect 3305 6951 3314 6971
rect 3344 6967 3407 6971
rect 3420 6967 3441 6973
rect 3344 6957 3398 6967
rect 3454 6951 3498 6985
rect 3503 6993 3532 7001
rect 3545 6993 3574 7058
rect 3873 7055 3907 7089
rect 3994 7067 4072 7089
rect 4106 7055 4120 7089
rect 4140 7083 4154 7123
rect 4506 7098 4668 7124
rect 4506 7097 4649 7098
rect 4506 7096 4536 7097
rect 4506 7055 4522 7096
rect 3585 6993 3600 7053
rect 3739 7025 3752 7053
rect 3697 7021 3833 7025
rect 3697 7013 3839 7021
rect 3697 7009 3752 7013
rect 3652 6993 3654 7009
rect 3686 6993 3688 7009
rect 3697 6993 3749 7009
rect 3773 6997 3839 7013
rect 3854 6997 3921 7052
rect 4007 7025 4038 7055
rect 4041 7039 4072 7055
rect 4041 7025 4158 7039
rect 3947 7021 3967 7025
rect 3979 7024 4001 7025
rect 4004 7024 4158 7025
rect 3941 7010 3967 7021
rect 3941 6997 3955 7010
rect 3970 7004 4158 7024
rect 3970 6997 4001 7004
rect 4007 6997 4158 7004
rect 3503 6978 3712 6993
rect 3503 6951 3697 6978
rect 3733 6951 3749 6993
rect 3752 6951 4158 6997
rect 1381 6926 1400 6938
rect 1447 6926 1454 6935
rect 1481 6926 1488 6935
rect 1493 6934 1523 6939
rect 1529 6934 1530 6939
rect 1493 6926 1530 6934
rect 1593 6936 1761 6941
rect 1593 6927 1663 6936
rect 1675 6935 1689 6936
rect 1711 6935 1761 6936
rect 1675 6933 1761 6935
rect 1770 6933 1830 6949
rect 1860 6941 4158 6951
rect 1860 6938 1889 6941
rect 1593 6926 1607 6927
rect 1616 6926 1655 6927
rect 1675 6926 1836 6933
rect 1110 6924 1836 6926
rect 1125 6920 1128 6924
rect 1153 6921 1163 6924
rect 1183 6923 1366 6924
rect 1142 6920 1163 6921
rect 960 6891 1183 6920
rect 968 6889 981 6891
rect 926 6884 981 6889
rect 994 6889 1183 6891
rect 1230 6904 1366 6923
rect 1230 6894 1351 6904
rect 1230 6889 1320 6894
rect 994 6885 1211 6889
rect 1241 6885 1286 6889
rect 994 6884 1286 6885
rect 926 6869 986 6884
rect 994 6874 1289 6884
rect 994 6873 1211 6874
rect 1025 6869 1122 6873
rect 1125 6869 1128 6873
rect 1142 6869 1211 6873
rect 1216 6873 1239 6874
rect 1241 6873 1289 6874
rect 1307 6873 1320 6889
rect 1216 6869 1351 6873
rect 926 6857 979 6869
rect 1013 6857 1211 6869
rect 965 6851 979 6857
rect 999 6853 1211 6857
rect 1217 6853 1351 6869
rect 1354 6863 1366 6904
rect 1381 6897 1400 6924
rect 1447 6901 1454 6924
rect 1478 6919 1530 6924
rect 1381 6884 1391 6897
rect 1478 6894 1523 6919
rect 1577 6918 1836 6924
rect 1860 6918 1874 6938
rect 1934 6936 4158 6941
rect 1936 6927 4158 6936
rect 1936 6926 2017 6927
rect 2023 6926 4158 6927
rect 1577 6899 1881 6918
rect 1934 6908 4158 6926
rect 1936 6907 4158 6908
rect 1478 6884 1490 6894
rect 1593 6891 1607 6899
rect 1616 6891 1881 6899
rect 1381 6873 1406 6884
rect 1478 6881 1505 6884
rect 1522 6881 1530 6887
rect 1478 6873 1530 6881
rect 1381 6872 1436 6873
rect 1443 6872 1532 6873
rect 1381 6869 1532 6872
rect 999 6851 1351 6853
rect 807 6846 1351 6851
rect 807 6831 1211 6846
rect 1217 6835 1351 6846
rect 1216 6831 1351 6835
rect 1406 6841 1436 6869
rect 1443 6841 1532 6869
rect 1406 6831 1532 6841
rect 1573 6831 1582 6891
rect 1593 6877 1881 6891
rect 1925 6899 4158 6907
rect 1925 6891 2003 6899
rect 1593 6857 1651 6877
rect 1675 6873 1881 6877
rect 1884 6873 1910 6881
rect 1925 6873 1944 6891
rect 1973 6884 2003 6891
rect 2006 6884 4158 6899
rect 1958 6877 4158 6884
rect 1958 6873 2018 6877
rect 2023 6873 4158 6877
rect 1675 6869 1914 6873
rect 1675 6861 1729 6869
rect 1744 6861 1784 6869
rect 1800 6861 1823 6869
rect 1850 6861 1857 6869
rect 1870 6861 1914 6869
rect 1593 6831 1645 6857
rect 1673 6831 1914 6861
rect 1925 6853 4158 6873
rect 9726 6858 9731 6892
rect 9726 6857 9765 6858
rect 1935 6837 4158 6853
rect 1935 6831 3347 6837
rect 807 6811 3347 6831
rect 3401 6819 3430 6837
rect 3545 6822 3554 6837
rect 3408 6811 3430 6819
rect 3442 6816 3534 6822
rect 3442 6811 3523 6816
rect 3622 6815 4158 6837
rect 807 6805 3344 6811
rect 817 6783 3344 6805
rect 859 6777 3344 6783
rect 859 6775 3347 6777
rect 3408 6775 3430 6777
rect 859 6750 3350 6775
rect 3442 6753 3512 6811
rect 3534 6777 3600 6796
rect 3622 6789 3642 6815
rect 3652 6793 3773 6811
rect 3820 6793 3962 6811
rect 3996 6793 4041 6811
rect 3534 6753 3566 6762
rect 552 6717 591 6749
rect 859 6748 3434 6750
rect 3442 6748 3566 6753
rect 859 6746 3566 6748
rect 859 6722 3350 6746
rect 3442 6743 3566 6746
rect 3354 6722 3384 6741
rect 859 6720 3406 6722
rect 3422 6720 3438 6725
rect 3442 6720 3534 6743
rect 859 6718 3552 6720
rect 859 6717 3350 6718
rect 921 6716 941 6717
rect 971 6716 1025 6717
rect 1008 6714 1025 6716
rect 796 6680 862 6700
rect 993 6699 1025 6714
rect 1038 6708 1062 6717
rect 1067 6708 1090 6717
rect 1008 6673 1013 6699
rect 1038 6680 1055 6708
rect 1103 6705 1137 6717
rect 1157 6705 1241 6717
rect 1103 6700 1171 6705
rect 1062 6680 1067 6700
rect 1103 6697 1198 6700
rect 1081 6691 1198 6697
rect 1267 6693 1276 6717
rect 1277 6695 1307 6717
rect 1242 6691 1267 6693
rect 1276 6691 1301 6693
rect 1081 6683 1264 6691
rect 1267 6683 1276 6691
rect 1346 6683 1347 6717
rect 1367 6709 1469 6717
rect 1367 6693 1432 6709
rect 1483 6707 1520 6717
rect 1533 6707 1565 6717
rect 1573 6707 1582 6717
rect 1611 6707 1646 6717
rect 1649 6707 1651 6717
rect 1441 6697 1507 6707
rect 1523 6703 1659 6707
rect 1081 6680 1276 6683
rect 1367 6681 1432 6691
rect 1441 6681 1519 6697
rect 1523 6692 1577 6703
rect 1607 6695 1659 6703
rect 1607 6692 1616 6695
rect 1646 6692 1659 6695
rect 1038 6675 1062 6680
rect 1039 6672 1062 6675
rect 1067 6672 1276 6680
rect 824 6652 862 6672
rect 1062 6652 1067 6672
rect 1081 6671 1276 6672
rect 1123 6663 1198 6671
rect 1205 6663 1276 6671
rect 1123 6659 1276 6663
rect 1124 6657 1276 6659
rect 1319 6657 1353 6681
rect 1367 6659 1519 6681
rect 1411 6657 1519 6659
rect 1533 6691 1577 6692
rect 1611 6691 1616 6692
rect 1649 6691 1651 6692
rect 1683 6691 1685 6717
rect 1725 6707 1857 6717
rect 1725 6705 1859 6707
rect 1711 6695 1859 6705
rect 1727 6692 1756 6695
rect 1765 6693 1859 6695
rect 1727 6691 1742 6692
rect 1533 6669 1616 6691
rect 1725 6685 1759 6691
rect 1533 6657 1577 6669
rect 1124 6653 1205 6657
rect 1124 6652 1242 6653
rect 1124 6641 1137 6652
rect 1176 6645 1242 6652
rect 1205 6641 1242 6645
rect 1441 6643 1543 6657
rect 1041 6639 1071 6641
rect 1205 6623 1276 6641
rect 1221 6619 1255 6623
rect 1313 6607 1347 6641
rect 1351 6627 1385 6643
rect 1423 6627 1543 6643
rect 1351 6623 1543 6627
rect 1351 6609 1545 6623
rect 1493 6597 1509 6609
rect 1517 6597 1545 6609
rect 1517 6593 1543 6597
rect 1559 6593 1583 6657
rect 1611 6623 1617 6657
rect 1649 6645 1651 6657
rect 1653 6623 1659 6685
rect 1725 6665 1763 6685
rect 1683 6627 1685 6657
rect 1691 6627 1697 6647
rect 1727 6638 1763 6665
rect 1777 6661 1859 6693
rect 1863 6691 1891 6717
rect 1973 6713 2003 6717
rect 2022 6713 2045 6717
rect 1893 6695 1912 6707
rect 1973 6695 1999 6713
rect 2017 6706 2045 6713
rect 2113 6707 2117 6717
rect 2135 6707 3350 6717
rect 2011 6695 2045 6706
rect 2071 6704 3350 6707
rect 2071 6697 2393 6704
rect 2053 6695 2393 6697
rect 1893 6692 2158 6695
rect 2162 6692 2177 6695
rect 2245 6692 2261 6695
rect 1893 6680 2099 6692
rect 1893 6669 2003 6680
rect 2011 6672 2099 6680
rect 1777 6645 1831 6661
rect 1914 6657 1927 6669
rect 1897 6649 1927 6657
rect 1777 6641 1807 6645
rect 1873 6641 1927 6649
rect 1931 6663 2003 6669
rect 2017 6663 2023 6672
rect 2027 6663 2099 6672
rect 1931 6657 2089 6663
rect 1931 6643 2071 6657
rect 2113 6652 2143 6692
rect 2260 6667 2261 6692
rect 2270 6671 2393 6695
rect 2417 6691 2422 6704
rect 2423 6695 2489 6704
rect 2423 6691 2492 6695
rect 2523 6691 2539 6704
rect 2562 6695 2564 6704
rect 2547 6691 2606 6695
rect 2631 6691 2708 6704
rect 2727 6695 2766 6704
rect 2751 6692 2766 6695
rect 2798 6691 3350 6704
rect 3354 6691 3384 6718
rect 3422 6707 3438 6718
rect 2291 6667 2393 6671
rect 2223 6657 2393 6667
rect 2423 6683 2523 6691
rect 2153 6652 2168 6657
rect 2260 6655 2261 6657
rect 2291 6655 2393 6657
rect 2301 6652 2331 6655
rect 2383 6652 2388 6655
rect 2417 6652 2422 6657
rect 2423 6655 2492 6683
rect 2547 6680 2688 6691
rect 2721 6681 3334 6691
rect 3388 6682 3406 6691
rect 3422 6682 3440 6707
rect 2562 6671 2688 6680
rect 2562 6655 2601 6671
rect 2631 6655 2688 6671
rect 2423 6652 2428 6655
rect 2490 6652 2492 6655
rect 2531 6652 2640 6655
rect 2658 6652 2688 6655
rect 2721 6657 2776 6676
rect 2798 6669 3334 6681
rect 2835 6657 3019 6669
rect 2721 6652 2742 6657
rect 2755 6652 2776 6657
rect 2873 6652 2945 6657
rect 2965 6652 3019 6657
rect 3073 6657 3207 6669
rect 3073 6652 3125 6657
rect 3133 6652 3212 6657
rect 3217 6652 3246 6657
rect 3442 6652 3534 6718
rect 1931 6641 2105 6643
rect 2113 6641 3650 6652
rect 1777 6638 3650 6641
rect 1727 6630 3650 6638
rect 1593 6593 1617 6623
rect 1683 6597 1723 6627
rect 1727 6626 3406 6630
rect 1727 6624 2346 6626
rect 2375 6624 2388 6626
rect 2658 6624 2673 6626
rect 2697 6624 2742 6626
rect 2755 6624 2776 6626
rect 2819 6624 3313 6626
rect 1727 6623 3622 6624
rect 1789 6597 1829 6623
rect 1832 6597 1849 6623
rect 1873 6619 1904 6623
rect 1931 6619 2037 6623
rect 1873 6597 1903 6619
rect 1927 6603 2037 6619
rect 2071 6609 2105 6623
rect 1927 6597 2003 6603
rect 2117 6602 3622 6623
rect 2117 6598 3434 6602
rect 1931 6595 2003 6597
rect 2275 6597 2341 6598
rect 2393 6597 2398 6598
rect 2520 6597 2522 6598
rect 2275 6593 2307 6597
rect 2309 6593 2341 6597
rect 2530 6593 2564 6598
rect 2598 6593 2640 6598
rect 2697 6597 2742 6598
rect 2721 6593 2742 6597
rect 2755 6593 2776 6598
rect 3125 6597 3155 6598
rect 3177 6597 3212 6598
rect 3183 6593 3212 6597
rect 3217 6597 3249 6598
rect 3217 6593 3246 6597
rect 1414 6575 1543 6593
rect 1649 6579 1723 6593
rect 1443 6571 1477 6575
rect 1645 6563 1723 6579
rect 1789 6587 1863 6593
rect 1789 6582 1873 6587
rect 1789 6563 1863 6582
rect 1645 6559 1697 6563
rect 1897 6561 2003 6593
rect 2052 6583 2068 6587
rect 2087 6583 2121 6593
rect 2037 6559 2153 6583
rect 2174 6582 2195 6587
rect 2249 6582 2301 6587
rect 2307 6565 2309 6593
rect 2375 6565 2422 6593
rect 2823 6589 3165 6593
rect 2873 6582 2891 6585
rect 2955 6582 2982 6585
rect 3123 6582 3170 6585
rect 3207 6582 3259 6585
rect 1645 6532 1663 6545
rect 2037 6532 2153 6549
rect 1414 6528 2826 6532
rect 1645 6525 1663 6528
rect 2037 6525 2153 6528
rect 1386 6500 2798 6504
rect 38 4296 1450 4300
rect 10 4268 1422 4272
rect 107 4207 205 4227
rect 255 4207 289 4229
rect 413 4207 492 4235
rect 496 4231 498 4245
rect 799 4231 802 4245
rect 496 4227 568 4231
rect 590 4227 676 4231
rect 496 4213 687 4227
rect 689 4213 802 4231
rect 936 4225 978 4231
rect 926 4223 978 4225
rect 829 4213 896 4223
rect 925 4213 978 4223
rect 268 4203 283 4207
rect 72 4189 102 4203
rect 257 4199 283 4203
rect 107 4189 205 4193
rect 72 4177 205 4189
rect 73 4175 205 4177
rect 241 4177 283 4199
rect 241 4175 285 4177
rect 78 4173 205 4175
rect 78 4159 180 4173
rect 215 4165 231 4175
rect 241 4169 279 4175
rect 269 4165 273 4169
rect 225 4163 231 4165
rect 117 4155 147 4159
rect 78 4125 90 4155
rect 112 4148 147 4155
rect 102 4118 147 4148
rect 102 4108 114 4118
rect 126 4111 146 4118
rect 126 4108 154 4111
rect 102 4096 154 4108
rect 23 4093 154 4096
rect 60 3999 72 4065
rect 126 4053 146 4093
rect 160 4036 180 4159
rect 217 4137 243 4163
rect 201 4036 206 4115
rect 156 4020 206 4036
rect 201 4019 206 4020
rect 217 4111 231 4137
rect 275 4115 279 4169
rect 309 4133 313 4207
rect 360 4157 374 4207
rect 496 4203 498 4213
rect 526 4207 602 4213
rect 623 4207 687 4213
rect 688 4203 689 4213
rect 447 4177 492 4201
rect 538 4177 540 4203
rect 560 4177 602 4193
rect 652 4191 653 4193
rect 619 4177 653 4191
rect 730 4177 731 4203
rect 799 4177 802 4213
rect 1025 4207 1137 4235
rect 1177 4213 1192 4231
rect 1198 4225 1264 4231
rect 1282 4229 1312 4231
rect 1267 4225 1312 4229
rect 1318 4225 1362 4231
rect 1198 4213 1362 4225
rect 1198 4207 1358 4213
rect 1392 4207 1422 4241
rect 1426 4235 1456 4275
rect 447 4173 653 4177
rect 394 4157 408 4173
rect 484 4169 653 4173
rect 484 4165 641 4169
rect 484 4162 513 4165
rect 217 4030 253 4111
rect 332 4110 460 4157
rect 484 4111 498 4162
rect 560 4131 641 4165
rect 568 4121 610 4131
rect 379 4105 460 4110
rect 481 4105 534 4111
rect 379 4093 454 4105
rect 484 4093 501 4105
rect 568 4093 646 4094
rect 379 4076 400 4093
rect 217 4024 231 4030
rect 235 4024 240 4030
rect 217 4009 246 4024
rect 273 4009 275 4047
rect 269 3999 275 4009
rect 307 3999 309 4013
rect 481 4011 500 4071
rect 515 4019 534 4077
rect 652 4029 653 4165
rect 676 4162 704 4177
rect 676 4108 689 4162
rect 762 4139 817 4177
rect 825 4139 827 4165
rect 873 4154 925 4169
rect 799 4131 817 4139
rect 873 4131 890 4154
rect 793 4108 890 4131
rect 676 4093 704 4108
rect 784 4105 890 4108
rect 784 4097 817 4105
rect 686 4079 687 4093
rect 676 4063 689 4079
rect 676 4049 724 4063
rect 730 4049 731 4093
rect 759 4071 846 4097
rect 687 4045 724 4049
rect 687 4037 732 4045
rect 758 4037 812 4063
rect 718 4029 732 4037
rect 413 3999 442 4011
rect 447 3999 481 4011
rect 515 3999 536 4019
rect 653 4003 732 4029
rect 758 4003 778 4029
rect 718 3999 732 4003
rect 765 3999 778 4003
rect 799 3999 812 4003
rect 813 3999 814 4071
rect 896 4056 925 4154
rect 1025 4139 1028 4207
rect 1041 4203 1056 4207
rect 1041 4201 1067 4203
rect 1123 4201 1144 4203
rect 1041 4177 1144 4201
rect 1198 4177 1204 4207
rect 1222 4181 1228 4203
rect 1232 4177 1324 4191
rect 1332 4177 1358 4207
rect 1059 4173 1137 4177
rect 1059 4139 1062 4173
rect 1093 4129 1094 4173
rect 1177 4162 1204 4177
rect 1227 4165 1374 4177
rect 1192 4133 1204 4162
rect 1232 4133 1238 4165
rect 1249 4162 1374 4165
rect 1192 4130 1198 4133
rect 1264 4131 1358 4162
rect 926 4114 1059 4121
rect 1093 4114 1114 4129
rect 1186 4121 1238 4130
rect 926 4105 1114 4114
rect 1017 4098 1022 4105
rect 944 4087 1025 4098
rect 1052 4087 1114 4105
rect 1173 4099 1238 4121
rect 1264 4115 1298 4131
rect 1312 4115 1318 4131
rect 926 4084 1114 4087
rect 926 4071 1059 4084
rect 881 4050 925 4056
rect 944 4051 1025 4071
rect 873 4043 976 4050
rect 981 4043 1025 4051
rect 1131 4043 1147 4053
rect 873 4041 1169 4043
rect 899 4038 1169 4041
rect 1173 4038 1181 4087
rect 1192 4086 1198 4099
rect 1220 4086 1238 4096
rect 1277 4086 1298 4115
rect 1332 4097 1358 4131
rect 1311 4086 1332 4097
rect 1188 4060 1332 4086
rect 1362 4063 1374 4162
rect 1460 4159 1517 4183
rect 1573 4159 1636 4183
rect 1697 4161 1749 4183
rect 1769 4170 1796 4183
rect 1769 4161 1811 4170
rect 1426 4125 1517 4149
rect 1552 4115 1561 4134
rect 1573 4115 1602 4149
rect 1768 4129 1775 4159
rect 1796 4155 1811 4161
rect 1836 4159 1937 4173
rect 2010 4159 2012 4193
rect 1796 4129 1822 4155
rect 1877 4139 1907 4155
rect 2044 4145 2046 4209
rect 2874 4200 4286 4204
rect 2846 4172 4258 4176
rect 1734 4114 1775 4129
rect 1345 4060 1374 4063
rect 1188 4039 1374 4060
rect 1207 4038 1215 4039
rect 0 3995 72 3999
rect 79 3995 368 3999
rect 0 3985 368 3995
rect 0 3961 72 3985
rect 79 3961 368 3985
rect 413 3987 604 3999
rect 627 3987 737 3999
rect 765 3995 884 3999
rect 413 3979 737 3987
rect 0 3957 368 3961
rect 418 3957 737 3979
rect 767 3979 884 3995
rect 899 3979 1220 4038
rect 767 3977 1220 3979
rect 1228 4021 1374 4039
rect 1521 4072 1577 4087
rect 1607 4081 1636 4091
rect 1717 4087 1725 4096
rect 1228 3999 1298 4021
rect 1311 4013 1374 4021
rect 1311 3999 1332 4013
rect 1345 3999 1374 4013
rect 1379 3999 1400 4029
rect 1459 4007 1519 4019
rect 1521 4018 1556 4072
rect 1561 4018 1577 4072
rect 1671 4065 1725 4087
rect 1749 4065 1775 4114
rect 1802 4065 1809 4129
rect 1870 4127 1937 4139
rect 1846 4125 1937 4127
rect 1846 4097 1873 4125
rect 1877 4117 1920 4125
rect 1938 4117 1968 4127
rect 1877 4097 1907 4117
rect 1937 4105 1968 4117
rect 1846 4065 1876 4097
rect 1938 4065 1968 4105
rect 2023 4097 2106 4129
rect 1521 4007 1577 4018
rect 1521 4003 1534 4007
rect 1546 4003 1577 4007
rect 1601 3999 1607 4059
rect 1671 4049 1775 4065
rect 1708 4015 1775 4049
rect 1667 3999 1670 4015
rect 1708 4003 1769 4015
rect 1799 4003 1877 4065
rect 1907 4015 1968 4065
rect 1973 4049 1983 4083
rect 2068 4075 2088 4077
rect 2119 4075 2122 4111
rect 2129 4097 2198 4129
rect 2267 4111 2398 4139
rect 2431 4123 2653 4135
rect 2491 4111 2653 4123
rect 2020 4045 2030 4049
rect 2034 4045 2054 4065
rect 2068 4045 2129 4075
rect 1983 4015 2129 4045
rect 1907 4003 2129 4015
rect 2153 4020 2156 4097
rect 2301 4077 2364 4105
rect 2572 4101 2593 4107
rect 2153 4011 2219 4020
rect 1708 3999 2224 4003
rect 1228 3989 1711 3999
rect 1228 3977 1270 3989
rect 743 3957 758 3973
rect 767 3957 1186 3977
rect 1198 3975 1225 3977
rect 1196 3957 1225 3975
rect 1277 3957 1711 3989
rect 1749 3957 2224 3999
rect -3 3947 2224 3957
rect 2267 3979 2287 4077
rect 2301 3979 2321 4077
rect 2428 4066 2446 4081
rect 2491 4077 2619 4101
rect 2671 4081 2701 4107
rect 2761 4077 2767 4101
rect 2796 4081 2807 4122
rect 2943 4111 3041 4131
rect 3091 4111 3125 4133
rect 3249 4111 3328 4139
rect 3332 4135 3334 4149
rect 3635 4135 3638 4149
rect 3332 4131 3404 4135
rect 3426 4131 3512 4135
rect 3332 4117 3523 4131
rect 3525 4117 3638 4135
rect 3772 4129 3814 4135
rect 3762 4127 3814 4129
rect 3665 4117 3732 4127
rect 3761 4117 3814 4127
rect 2510 4066 2530 4077
rect 2603 4067 2623 4077
rect 2428 4051 2431 4066
rect 2420 4048 2470 4051
rect 2510 4048 2515 4066
rect 2551 4048 2554 4067
rect 2585 4048 2588 4067
rect 2613 4049 2623 4067
rect 2727 4049 2733 4077
rect 2761 4067 2795 4077
rect 2761 4051 2767 4067
rect 2814 4051 2819 4111
rect 2602 4048 2623 4049
rect 2420 4019 2643 4048
rect 2428 4017 2441 4019
rect 2386 4012 2441 4017
rect 2454 4017 2643 4019
rect 2701 4017 2733 4049
rect 2848 4025 2853 4111
rect 3104 4107 3119 4111
rect 2908 4093 2938 4107
rect 3093 4103 3119 4107
rect 2943 4093 3041 4097
rect 2908 4081 3041 4093
rect 2909 4079 3041 4081
rect 3077 4081 3119 4103
rect 3077 4079 3121 4081
rect 2914 4077 3041 4079
rect 2914 4063 3016 4077
rect 3051 4069 3067 4079
rect 3077 4073 3115 4079
rect 3105 4069 3109 4073
rect 3061 4067 3067 4069
rect 2953 4059 2983 4063
rect 2914 4029 2926 4059
rect 2948 4052 2983 4059
rect 2938 4022 2983 4052
rect 2386 3997 2446 4012
rect 2454 4001 2671 4017
rect 2701 4012 2731 4017
rect 2938 4012 2950 4022
rect 2962 4015 2982 4022
rect 2962 4012 2990 4015
rect 2485 3997 2582 4001
rect 2585 3997 2588 4001
rect 2602 3997 2671 4001
rect 2677 3997 2699 4011
rect 2701 3997 2746 4012
rect 2938 4000 2990 4012
rect 2859 3997 2990 4000
rect 2386 3985 2439 3997
rect 2473 3985 2875 3997
rect 2425 3979 2439 3985
rect 2459 3979 2875 3985
rect -3 3941 2266 3947
rect 117 3931 144 3941
rect 157 3931 189 3941
rect 201 3931 206 3941
rect 235 3931 240 3941
rect 65 3927 117 3931
rect 147 3927 240 3931
rect 65 3917 201 3927
rect 65 3893 143 3917
rect 147 3916 201 3917
rect 157 3893 201 3916
rect 235 3919 240 3927
rect 65 3881 207 3893
rect 65 3855 167 3881
rect 47 3851 167 3855
rect 4 3847 167 3851
rect 4 3833 169 3847
rect 117 3821 133 3833
rect 141 3821 169 3833
rect 141 3817 167 3821
rect 183 3817 207 3881
rect 235 3847 241 3919
rect 273 3869 275 3941
rect 277 3847 283 3909
rect 307 3851 309 3941
rect 453 3931 486 3941
rect 353 3929 483 3931
rect 353 3916 368 3929
rect 373 3919 483 3929
rect 389 3917 483 3919
rect 315 3851 321 3871
rect 351 3862 387 3909
rect 401 3885 483 3917
rect 487 3895 515 3941
rect 743 3931 758 3941
rect 777 3931 812 3939
rect 517 3919 536 3931
rect 695 3921 812 3931
rect 677 3919 812 3921
rect 846 3931 944 3941
rect 967 3931 1017 3941
rect 846 3919 1017 3931
rect 517 3904 647 3919
rect 517 3893 627 3904
rect 401 3869 455 3885
rect 521 3873 551 3893
rect 401 3865 431 3869
rect 497 3865 551 3873
rect 555 3887 627 3893
rect 641 3887 647 3904
rect 651 3916 792 3919
rect 869 3916 885 3919
rect 651 3887 723 3916
rect 555 3865 695 3887
rect 737 3865 767 3916
rect 777 3865 792 3916
rect 884 3879 885 3916
rect 894 3895 1017 3919
rect 915 3879 1017 3895
rect 925 3865 955 3879
rect 401 3862 970 3865
rect 217 3817 241 3847
rect 307 3821 347 3851
rect 351 3847 970 3862
rect 1007 3851 1012 3879
rect 1041 3855 1046 3941
rect 1047 3919 1113 3941
rect 1186 3919 1188 3941
rect 1277 3931 1298 3941
rect 1311 3931 1351 3941
rect 1379 3939 1400 3941
rect 1271 3929 1332 3931
rect 1047 3879 1116 3919
rect 1171 3907 1230 3919
rect 1255 3907 1332 3929
rect 1171 3904 1312 3907
rect 1186 3895 1312 3904
rect 1186 3879 1225 3895
rect 1255 3879 1312 3895
rect 1047 3857 1052 3879
rect 1114 3857 1116 3879
rect 1061 3855 1095 3857
rect 1155 3851 1264 3879
rect 1282 3857 1312 3879
rect 1345 3857 1366 3885
rect 413 3821 453 3847
rect 456 3821 473 3847
rect 497 3843 528 3847
rect 555 3843 661 3847
rect 497 3821 527 3843
rect 551 3827 661 3843
rect 695 3833 729 3847
rect 777 3827 792 3847
rect 551 3821 627 3827
rect 925 3823 955 3847
rect 999 3823 1012 3851
rect 1282 3847 1297 3857
rect 555 3819 627 3821
rect 899 3821 965 3823
rect 1017 3821 1022 3847
rect 1144 3821 1146 3847
rect 1228 3845 1255 3847
rect 899 3817 931 3821
rect 933 3817 965 3821
rect 1154 3817 1188 3845
rect 1222 3817 1264 3845
rect 1321 3821 1366 3857
rect 1345 3817 1366 3821
rect 1379 3817 1400 3900
rect 1422 3893 2266 3941
rect 2267 3933 2875 3979
rect 2277 3911 2875 3933
rect 1498 3881 1608 3893
rect 1520 3862 1608 3881
rect 1505 3851 1622 3862
rect 1627 3859 1635 3893
rect 1639 3881 1643 3893
rect 1477 3847 1622 3851
rect 1661 3851 1669 3893
rect 1697 3881 1846 3893
rect 1677 3851 1681 3881
rect 1697 3869 1755 3881
rect 1697 3863 1749 3869
rect 1761 3863 1846 3881
rect 1853 3863 1870 3893
rect 1876 3863 1907 3893
rect 2012 3863 2266 3893
rect 1697 3858 2266 3863
rect 2319 3903 2875 3911
rect 2896 3903 2908 3969
rect 2962 3957 2982 3997
rect 2996 3940 3016 4063
rect 3053 4041 3079 4067
rect 3037 3940 3042 4019
rect 2992 3924 3042 3940
rect 3037 3923 3042 3924
rect 3053 4015 3067 4041
rect 3111 4019 3115 4073
rect 3145 4037 3149 4111
rect 3196 4061 3210 4111
rect 3332 4107 3334 4117
rect 3362 4111 3438 4117
rect 3459 4111 3523 4117
rect 3524 4107 3525 4117
rect 3283 4081 3328 4105
rect 3374 4081 3376 4107
rect 3396 4081 3438 4097
rect 3488 4095 3489 4097
rect 3455 4081 3489 4095
rect 3566 4081 3567 4107
rect 3635 4081 3638 4117
rect 3861 4111 3973 4139
rect 4013 4117 4028 4135
rect 4034 4129 4100 4135
rect 4118 4133 4148 4135
rect 4103 4129 4148 4133
rect 4154 4129 4198 4135
rect 4034 4117 4198 4129
rect 4034 4111 4194 4117
rect 4228 4111 4258 4145
rect 4262 4139 4292 4179
rect 3283 4077 3489 4081
rect 3230 4061 3244 4077
rect 3320 4073 3489 4077
rect 3320 4069 3477 4073
rect 3320 4066 3349 4069
rect 3053 3934 3089 4015
rect 3168 4014 3296 4061
rect 3320 4015 3334 4066
rect 3396 4035 3477 4069
rect 3404 4025 3446 4035
rect 3215 4009 3296 4014
rect 3317 4009 3370 4015
rect 3215 3997 3290 4009
rect 3320 3997 3337 4009
rect 3404 3997 3482 3998
rect 3215 3980 3236 3997
rect 3053 3928 3067 3934
rect 3071 3928 3076 3934
rect 3053 3913 3082 3928
rect 3109 3913 3111 3951
rect 3105 3903 3111 3913
rect 3143 3903 3145 3917
rect 3317 3915 3336 3975
rect 3351 3923 3370 3981
rect 3488 3933 3489 4069
rect 3512 4066 3540 4081
rect 3512 4012 3525 4066
rect 3598 4043 3653 4081
rect 3661 4043 3663 4069
rect 3709 4058 3761 4073
rect 3635 4035 3653 4043
rect 3709 4035 3726 4058
rect 3629 4012 3726 4035
rect 3512 3997 3540 4012
rect 3620 4009 3726 4012
rect 3620 4001 3653 4009
rect 3522 3983 3523 3997
rect 3512 3967 3525 3983
rect 3512 3953 3560 3967
rect 3566 3953 3567 3997
rect 3595 3975 3682 4001
rect 3523 3949 3560 3953
rect 3523 3941 3568 3949
rect 3594 3941 3648 3967
rect 3554 3933 3568 3941
rect 3249 3903 3278 3915
rect 3283 3903 3317 3915
rect 3351 3903 3372 3923
rect 3489 3907 3568 3933
rect 3594 3907 3614 3933
rect 3554 3903 3568 3907
rect 3601 3903 3614 3907
rect 3635 3903 3648 3907
rect 3649 3903 3650 3975
rect 3732 3960 3761 4058
rect 3861 4043 3864 4111
rect 3877 4107 3892 4111
rect 3877 4105 3903 4107
rect 3959 4105 3980 4107
rect 3877 4081 3980 4105
rect 4034 4081 4040 4111
rect 4058 4085 4064 4107
rect 4068 4081 4160 4095
rect 4168 4081 4194 4111
rect 4585 4087 4615 4101
rect 3895 4077 3973 4081
rect 3895 4043 3898 4077
rect 3929 4033 3930 4077
rect 4013 4066 4040 4081
rect 4063 4069 4210 4081
rect 4028 4037 4040 4066
rect 4068 4037 4074 4069
rect 4085 4066 4210 4069
rect 4028 4034 4034 4037
rect 4100 4035 4194 4066
rect 3762 4018 3895 4025
rect 3929 4018 3950 4033
rect 4022 4025 4074 4034
rect 3762 4009 3950 4018
rect 3853 4002 3858 4009
rect 3780 3991 3861 4002
rect 3888 3991 3950 4009
rect 4009 4003 4074 4025
rect 4100 4019 4134 4035
rect 4148 4019 4154 4035
rect 3762 3988 3950 3991
rect 3762 3975 3895 3988
rect 3717 3954 3761 3960
rect 3780 3955 3861 3975
rect 3709 3947 3812 3954
rect 3817 3947 3861 3955
rect 3967 3947 3983 3957
rect 3709 3945 4005 3947
rect 3735 3942 4005 3945
rect 4009 3942 4017 3991
rect 4028 3990 4034 4003
rect 4056 3990 4074 4000
rect 4113 3990 4134 4019
rect 4168 4001 4194 4035
rect 4147 3990 4168 4001
rect 4024 3964 4168 3990
rect 4198 3967 4210 4066
rect 4296 4063 4322 4087
rect 4375 4063 4472 4087
rect 4533 4065 4632 4087
rect 4427 4059 4432 4063
rect 4262 4029 4322 4053
rect 4375 4033 4443 4053
rect 4469 4033 4474 4059
rect 4181 3964 4210 3967
rect 4024 3943 4210 3964
rect 4043 3942 4051 3943
rect 2319 3899 2908 3903
rect 2915 3899 3204 3903
rect 2319 3889 3204 3899
rect 2319 3865 2908 3889
rect 2915 3865 3204 3889
rect 3249 3891 3440 3903
rect 3463 3891 3573 3903
rect 3601 3899 3720 3903
rect 3249 3883 3573 3891
rect 2319 3861 3204 3865
rect 3254 3861 3573 3883
rect 3603 3883 3720 3899
rect 3735 3883 4056 3942
rect 3603 3881 4056 3883
rect 4064 3925 4210 3943
rect 4333 4018 4351 4033
rect 4363 4029 4469 4033
rect 4363 4018 4385 4029
rect 4333 3992 4336 4018
rect 4378 4003 4385 4018
rect 4388 4019 4469 4029
rect 4388 4017 4404 4019
rect 4406 4018 4447 4019
rect 4406 4017 4437 4018
rect 4333 3961 4341 3992
rect 4064 3903 4134 3925
rect 4147 3917 4210 3925
rect 4147 3903 4168 3917
rect 4181 3903 4210 3917
rect 4215 3903 4236 3933
rect 4333 3919 4355 3961
rect 4375 3919 4403 3985
rect 4333 3911 4403 3919
rect 4322 3903 4355 3911
rect 4064 3893 4374 3903
rect 4064 3881 4106 3893
rect 3579 3861 3594 3877
rect 3603 3861 4022 3881
rect 4034 3879 4061 3881
rect 4032 3861 4061 3879
rect 4113 3861 4374 3893
rect 4375 3861 4403 3911
rect 4409 3861 4437 4017
rect 4475 3969 4506 4063
rect 4509 4000 4540 4063
rect 4585 4033 4615 4065
rect 4719 4063 4756 4077
rect 4643 4059 4672 4063
rect 4637 4033 4672 4059
rect 4583 4021 4630 4033
rect 4583 4018 4627 4021
rect 4585 4000 4615 4018
rect 4509 3987 4627 4000
rect 4507 3969 4635 3987
rect 4643 3969 4672 4033
rect 4677 4033 4706 4063
rect 4677 4031 4709 4033
rect 4677 3984 4712 4031
rect 4719 4029 4773 4043
rect 4722 4009 4745 4029
rect 4677 3971 4719 3984
rect 4682 3969 4719 3971
rect 4507 3953 4637 3969
rect 4475 3903 4506 3919
rect 4509 3915 4540 3919
rect 4509 3903 4543 3915
rect 4544 3903 4553 3953
rect 4554 3919 4637 3953
rect 4643 3949 4719 3969
rect 4643 3937 4794 3949
rect 4583 3907 4637 3919
rect 4667 3907 4794 3937
rect 5082 3917 5102 3949
rect 4583 3903 4794 3907
rect 4541 3869 4577 3881
rect 4585 3861 4794 3903
rect 1697 3851 2224 3858
rect 1661 3847 2224 3851
rect 1520 3831 1542 3847
rect 1749 3835 1789 3847
rect 1749 3831 1769 3835
rect 1819 3817 1836 3847
rect 1853 3817 1870 3847
rect 1877 3821 1907 3831
rect 1938 3821 1949 3847
rect 2012 3845 2224 3847
rect 2072 3821 2094 3845
rect 2122 3817 2138 3845
rect 2156 3839 2178 3845
rect 2156 3836 2206 3839
rect 2156 3817 2217 3836
rect 2253 3828 2280 3851
rect 2319 3845 4794 3861
rect 2381 3844 2401 3845
rect 2431 3844 2485 3845
rect 2468 3842 2485 3844
rect 2453 3828 2485 3842
rect 2498 3828 2515 3845
rect 2563 3833 2597 3845
rect 2617 3833 2701 3845
rect 2953 3835 2980 3845
rect 2993 3835 3025 3845
rect 3037 3835 3042 3845
rect 3071 3835 3076 3845
rect 2563 3828 2631 3833
rect 2901 3831 2953 3835
rect 2983 3831 3076 3835
rect 38 3799 167 3817
rect 273 3803 347 3817
rect 67 3795 101 3799
rect 269 3787 347 3803
rect 413 3811 487 3817
rect 413 3806 497 3811
rect 413 3787 487 3806
rect 269 3783 321 3787
rect 521 3785 627 3817
rect 676 3807 692 3811
rect 711 3807 745 3817
rect 661 3783 777 3807
rect 798 3806 819 3811
rect 873 3806 925 3811
rect 931 3789 933 3817
rect 999 3789 1046 3817
rect 1447 3813 1757 3817
rect 1734 3806 1769 3809
rect 1831 3806 1877 3809
rect 1923 3806 1983 3809
rect 2172 3805 2217 3817
rect 2183 3783 2217 3805
rect 2219 3783 2246 3817
rect 2253 3808 2527 3828
rect 2563 3825 2864 3828
rect 2541 3808 2864 3825
rect 2901 3821 3037 3831
rect 269 3756 287 3769
rect 661 3756 777 3773
rect 38 3752 1450 3756
rect 269 3749 287 3752
rect 661 3749 777 3752
rect 2253 3749 2280 3808
rect 2468 3801 2473 3808
rect 2498 3803 2515 3808
rect 2541 3807 2727 3808
rect 2539 3805 2727 3807
rect 2541 3803 2727 3805
rect 2540 3801 2724 3803
rect 2541 3800 2724 3801
rect 2736 3800 2761 3808
rect 2284 3780 2527 3800
rect 2541 3799 2836 3800
rect 2583 3787 2836 3799
rect 2584 3780 2836 3787
rect 2901 3797 2979 3821
rect 2983 3820 3037 3821
rect 2993 3797 3037 3820
rect 3071 3823 3076 3831
rect 2901 3785 3043 3797
rect 2584 3769 2597 3780
rect 2636 3773 2702 3780
rect 2665 3769 2702 3773
rect 2736 3769 2761 3780
rect 2501 3767 2531 3769
rect 2773 3735 2807 3769
rect 2811 3755 2845 3771
rect 2901 3759 3003 3785
rect 2883 3755 3003 3759
rect 2811 3751 3003 3755
rect 2811 3737 3005 3751
rect 10 3724 1422 3728
rect 2953 3725 2969 3737
rect 2977 3725 3005 3737
rect 2977 3721 3003 3725
rect 3019 3721 3043 3785
rect 3071 3751 3077 3823
rect 3109 3773 3111 3845
rect 3113 3751 3119 3813
rect 3143 3755 3145 3845
rect 3289 3835 3322 3845
rect 3189 3833 3319 3835
rect 3189 3820 3204 3833
rect 3209 3823 3319 3833
rect 3225 3821 3319 3823
rect 3151 3755 3157 3775
rect 3187 3766 3223 3813
rect 3237 3789 3319 3821
rect 3323 3799 3351 3845
rect 3579 3835 3594 3845
rect 3613 3835 3648 3843
rect 3353 3823 3372 3835
rect 3531 3825 3648 3835
rect 3513 3823 3648 3825
rect 3682 3835 3780 3845
rect 3803 3835 3853 3845
rect 3682 3823 3853 3835
rect 3353 3808 3483 3823
rect 3353 3797 3463 3808
rect 3237 3773 3291 3789
rect 3357 3777 3387 3797
rect 3237 3769 3267 3773
rect 3333 3769 3387 3777
rect 3391 3791 3463 3797
rect 3477 3791 3483 3808
rect 3487 3820 3628 3823
rect 3705 3820 3721 3823
rect 3487 3791 3559 3820
rect 3391 3769 3531 3791
rect 3573 3769 3603 3820
rect 3613 3769 3628 3820
rect 3720 3783 3721 3820
rect 3730 3799 3853 3823
rect 3751 3783 3853 3799
rect 3761 3769 3791 3783
rect 3237 3766 3806 3769
rect 3053 3721 3077 3751
rect 3143 3725 3183 3755
rect 3187 3751 3806 3766
rect 3843 3755 3848 3783
rect 3877 3759 3882 3845
rect 3883 3823 3949 3845
rect 4022 3823 4024 3845
rect 4113 3835 4134 3845
rect 4147 3835 4187 3845
rect 4215 3843 4236 3845
rect 4107 3833 4168 3835
rect 3883 3783 3952 3823
rect 4007 3811 4066 3823
rect 4091 3811 4168 3833
rect 4007 3808 4148 3811
rect 4022 3799 4148 3808
rect 4022 3783 4061 3799
rect 4091 3783 4148 3799
rect 3883 3761 3888 3783
rect 3950 3761 3952 3783
rect 3897 3759 3931 3761
rect 3991 3755 4100 3783
rect 4118 3761 4148 3783
rect 4181 3761 4202 3789
rect 3249 3725 3289 3751
rect 3292 3725 3309 3751
rect 3333 3747 3364 3751
rect 3391 3747 3497 3751
rect 3333 3725 3363 3747
rect 3387 3731 3497 3747
rect 3531 3737 3565 3751
rect 3613 3731 3628 3751
rect 3387 3725 3463 3731
rect 3761 3727 3791 3751
rect 3835 3727 3848 3755
rect 4118 3751 4133 3761
rect 3391 3723 3463 3725
rect 3735 3725 3801 3727
rect 3853 3725 3858 3751
rect 3980 3725 3982 3751
rect 4064 3749 4091 3751
rect 3735 3721 3767 3725
rect 3769 3721 3801 3725
rect 3990 3721 4024 3749
rect 4058 3721 4100 3749
rect 4157 3725 4202 3761
rect 4181 3721 4202 3725
rect 4215 3721 4236 3804
rect 4258 3797 4794 3845
rect 4295 3785 4479 3797
rect 4333 3767 4405 3785
rect 4425 3767 4479 3785
rect 4279 3755 4479 3767
rect 4533 3785 4672 3797
rect 4533 3767 4585 3785
rect 4593 3767 4672 3785
rect 4677 3767 4706 3797
rect 4533 3755 4773 3767
rect 4279 3751 4773 3755
rect 4643 3735 4672 3751
rect 4585 3725 4615 3735
rect 4637 3725 4672 3735
rect 4643 3721 4672 3725
rect 4677 3725 4709 3751
rect 4677 3721 4706 3725
rect 2874 3703 3003 3721
rect 3109 3707 3183 3721
rect 2903 3699 2937 3703
rect 3105 3691 3183 3707
rect 3249 3715 3323 3721
rect 3249 3710 3333 3715
rect 3249 3691 3323 3710
rect 3105 3687 3157 3691
rect 3357 3689 3463 3721
rect 3512 3711 3528 3715
rect 3547 3711 3581 3721
rect 3497 3687 3613 3711
rect 3634 3710 3655 3715
rect 3709 3710 3761 3715
rect 3767 3693 3769 3721
rect 3835 3693 3882 3721
rect 4283 3717 4625 3721
rect 4333 3710 4351 3713
rect 4415 3710 4442 3713
rect 4583 3710 4630 3713
rect 4667 3710 4719 3713
rect 3105 3660 3123 3673
rect 3497 3660 3613 3677
rect 2874 3656 4286 3660
rect 3105 3653 3123 3656
rect 3497 3653 3613 3656
rect 2846 3628 4258 3632
rect 12648 3562 12852 3564
rect 1220 3408 1486 3412
rect 1536 3408 2620 3412
rect 1220 3380 1486 3384
rect 1494 3382 1530 3392
rect 1536 3382 2592 3384
rect 1494 3380 2592 3382
rect 1456 3341 1459 3353
rect 1494 3348 1551 3380
rect 2562 3364 2592 3366
rect 2596 3364 2626 3400
rect 2750 3394 2752 3397
rect 2716 3360 2718 3364
rect 2750 3363 2799 3394
rect 1277 3319 1375 3339
rect 1425 3319 1459 3341
rect 1517 3319 1551 3348
rect 1583 3319 1662 3347
rect 1666 3343 1668 3357
rect 1969 3343 1972 3357
rect 1666 3339 1738 3343
rect 1760 3339 1846 3343
rect 1666 3325 1857 3339
rect 1859 3325 1972 3343
rect 2106 3337 2148 3343
rect 2096 3335 2148 3337
rect 1999 3325 2066 3335
rect 2095 3325 2148 3335
rect 1438 3315 1453 3319
rect 1242 3301 1272 3315
rect 1427 3311 1453 3315
rect 1277 3301 1375 3305
rect 1242 3289 1375 3301
rect 1243 3287 1375 3289
rect 1411 3289 1453 3311
rect 1411 3287 1455 3289
rect 1248 3285 1375 3287
rect 1248 3271 1350 3285
rect 1385 3277 1401 3287
rect 1411 3281 1449 3287
rect 1439 3277 1443 3281
rect 1395 3275 1401 3277
rect 1287 3267 1317 3271
rect 1248 3237 1260 3267
rect 1282 3260 1317 3267
rect 1272 3230 1317 3260
rect 1272 3220 1284 3230
rect 1296 3223 1316 3230
rect 1296 3220 1324 3223
rect 1272 3208 1324 3220
rect 1193 3205 1324 3208
rect 1230 3111 1242 3177
rect 1296 3165 1316 3205
rect 1330 3148 1350 3271
rect 1387 3249 1413 3275
rect 1371 3148 1376 3227
rect 1326 3132 1376 3148
rect 1371 3131 1376 3132
rect 1387 3223 1401 3249
rect 1445 3227 1449 3281
rect 1479 3245 1483 3319
rect 1530 3269 1544 3319
rect 1666 3315 1668 3325
rect 1696 3319 1772 3325
rect 1793 3319 1857 3325
rect 1858 3315 1859 3325
rect 1617 3289 1662 3313
rect 1708 3289 1710 3315
rect 1730 3289 1772 3305
rect 1822 3303 1823 3305
rect 1789 3289 1823 3303
rect 1900 3289 1901 3315
rect 1969 3289 1972 3325
rect 2195 3319 2307 3347
rect 2347 3325 2362 3343
rect 2368 3337 2434 3343
rect 2452 3341 2482 3343
rect 2437 3337 2482 3341
rect 2488 3337 2532 3343
rect 2368 3325 2532 3337
rect 2688 3326 2765 3360
rect 2731 3325 2765 3326
rect 2368 3319 2528 3325
rect 1617 3285 1823 3289
rect 1564 3269 1578 3285
rect 1654 3281 1823 3285
rect 1654 3277 1811 3281
rect 1654 3274 1683 3277
rect 1387 3142 1423 3223
rect 1502 3222 1630 3269
rect 1654 3223 1668 3274
rect 1730 3243 1811 3277
rect 1738 3233 1780 3243
rect 1549 3217 1630 3222
rect 1651 3217 1704 3223
rect 1549 3205 1624 3217
rect 1654 3205 1671 3217
rect 1738 3205 1816 3206
rect 1549 3188 1570 3205
rect 1387 3136 1401 3142
rect 1405 3136 1410 3142
rect 1387 3121 1416 3136
rect 1443 3121 1445 3159
rect 1439 3111 1445 3121
rect 1477 3111 1479 3125
rect 1651 3123 1670 3183
rect 1685 3131 1704 3189
rect 1822 3141 1823 3277
rect 1846 3274 1874 3289
rect 1846 3220 1859 3274
rect 1932 3251 1987 3289
rect 1995 3251 1997 3277
rect 2043 3266 2095 3281
rect 1969 3243 1987 3251
rect 2043 3243 2060 3266
rect 1963 3220 2060 3243
rect 1846 3205 1874 3220
rect 1954 3217 2060 3220
rect 1954 3209 1987 3217
rect 1856 3191 1857 3205
rect 1846 3175 1859 3191
rect 1846 3161 1894 3175
rect 1900 3161 1901 3205
rect 1929 3183 2016 3209
rect 1857 3157 1894 3161
rect 1857 3149 1902 3157
rect 1928 3149 1982 3175
rect 1888 3141 1902 3149
rect 1583 3111 1612 3123
rect 1617 3111 1651 3123
rect 1685 3111 1706 3131
rect 1823 3115 1902 3141
rect 1928 3115 1948 3141
rect 1888 3111 1902 3115
rect 1935 3111 1948 3115
rect 1969 3111 1982 3115
rect 1983 3111 1984 3183
rect 2066 3168 2095 3266
rect 2195 3251 2198 3319
rect 2211 3315 2226 3319
rect 2211 3313 2237 3315
rect 2293 3313 2314 3315
rect 2211 3289 2314 3313
rect 2368 3289 2374 3319
rect 2392 3293 2398 3315
rect 2402 3289 2494 3303
rect 2502 3289 2528 3319
rect 2229 3285 2307 3289
rect 2229 3251 2232 3285
rect 2263 3241 2264 3285
rect 2347 3274 2374 3289
rect 2397 3277 2544 3289
rect 2362 3245 2374 3274
rect 2402 3245 2408 3277
rect 2419 3274 2544 3277
rect 2362 3242 2368 3245
rect 2434 3243 2528 3274
rect 2096 3226 2229 3233
rect 2263 3226 2284 3241
rect 2356 3233 2408 3242
rect 2096 3217 2284 3226
rect 2187 3210 2192 3217
rect 2114 3199 2195 3210
rect 2222 3199 2284 3217
rect 2343 3211 2408 3233
rect 2434 3227 2468 3243
rect 2482 3227 2488 3243
rect 2096 3196 2284 3199
rect 2096 3183 2229 3196
rect 2051 3162 2095 3168
rect 2114 3163 2195 3183
rect 2043 3155 2146 3162
rect 2151 3155 2195 3163
rect 2301 3155 2317 3165
rect 2043 3153 2339 3155
rect 2069 3150 2339 3153
rect 2343 3150 2351 3199
rect 2362 3198 2368 3211
rect 2390 3198 2408 3208
rect 2447 3198 2468 3227
rect 2502 3209 2528 3243
rect 2481 3198 2502 3209
rect 2358 3172 2502 3198
rect 2532 3175 2544 3274
rect 2515 3172 2544 3175
rect 2731 3288 2754 3325
rect 2731 3172 2765 3288
rect 2358 3151 2544 3172
rect 2377 3150 2385 3151
rect 1167 3107 1242 3111
rect 1249 3107 1538 3111
rect 1167 3097 1538 3107
rect 1167 3073 1242 3097
rect 1249 3073 1538 3097
rect 1583 3099 1774 3111
rect 1797 3099 1907 3111
rect 1935 3107 2054 3111
rect 1583 3091 1907 3099
rect 1167 3069 1538 3073
rect 1588 3069 1907 3091
rect 1937 3091 2054 3107
rect 2069 3091 2390 3150
rect 1937 3089 2390 3091
rect 2398 3133 2544 3151
rect 2688 3169 2765 3172
rect 2398 3111 2468 3133
rect 2481 3125 2544 3133
rect 2481 3111 2502 3125
rect 2515 3111 2544 3125
rect 2549 3111 2570 3141
rect 2688 3138 2717 3169
rect 2731 3149 2765 3169
rect 2720 3138 2765 3149
rect 2771 3111 2799 3171
rect 3038 3118 3080 3128
rect 3040 3114 3080 3118
rect 2398 3101 2828 3111
rect 2398 3089 2440 3101
rect 1913 3069 1928 3085
rect 1937 3069 2356 3089
rect 2368 3087 2395 3089
rect 2366 3069 2395 3087
rect 2447 3088 2828 3101
rect 3010 3090 3052 3100
rect 2447 3069 2826 3088
rect 3012 3086 3052 3090
rect 1167 3064 2826 3069
rect 1167 3053 2630 3064
rect 1287 3043 1314 3053
rect 1327 3043 1359 3053
rect 1371 3043 1376 3053
rect 1405 3043 1410 3053
rect 1235 3039 1287 3043
rect 1317 3039 1410 3043
rect 1235 3029 1371 3039
rect 1235 3005 1313 3029
rect 1317 3028 1371 3029
rect 1327 3005 1371 3028
rect 1405 3031 1410 3039
rect 1235 2993 1377 3005
rect 1235 2967 1337 2993
rect 1217 2963 1337 2967
rect 1174 2959 1337 2963
rect 1174 2945 1339 2959
rect 1287 2933 1303 2945
rect 1311 2933 1339 2945
rect 1311 2929 1337 2933
rect 1353 2929 1377 2993
rect 1405 2959 1411 3031
rect 1443 2981 1445 3053
rect 1447 2959 1453 3021
rect 1477 2963 1479 3053
rect 1623 3043 1656 3053
rect 1523 3041 1653 3043
rect 1523 3028 1538 3041
rect 1543 3031 1653 3041
rect 1559 3029 1653 3031
rect 1485 2963 1491 2983
rect 1521 2974 1557 3021
rect 1571 2997 1653 3029
rect 1657 3007 1685 3053
rect 1913 3043 1928 3053
rect 1947 3043 1982 3051
rect 1687 3031 1706 3043
rect 1865 3033 1982 3043
rect 1847 3031 1982 3033
rect 2016 3043 2114 3053
rect 2137 3043 2187 3053
rect 2016 3031 2187 3043
rect 1687 3016 1817 3031
rect 1687 3005 1797 3016
rect 1571 2981 1625 2997
rect 1691 2985 1721 3005
rect 1571 2977 1601 2981
rect 1667 2977 1721 2985
rect 1725 2999 1797 3005
rect 1811 2999 1817 3016
rect 1821 3028 1962 3031
rect 2039 3028 2055 3031
rect 1821 2999 1893 3028
rect 1725 2977 1865 2999
rect 1907 2977 1937 3028
rect 1947 2977 1962 3028
rect 2054 2991 2055 3028
rect 2064 3007 2187 3031
rect 2085 2991 2187 3007
rect 2211 3052 2288 3053
rect 2211 3040 2290 3052
rect 2095 2977 2125 2991
rect 1571 2974 2140 2977
rect 1387 2929 1411 2959
rect 1477 2933 1517 2963
rect 1521 2959 2140 2974
rect 2177 2963 2182 2991
rect 2211 2967 2216 3040
rect 2217 3031 2283 3040
rect 2356 3031 2358 3053
rect 2447 3043 2468 3053
rect 2481 3043 2521 3053
rect 2549 3051 2570 3053
rect 2441 3041 2502 3043
rect 2217 2991 2286 3031
rect 2341 3019 2400 3031
rect 2425 3019 2502 3041
rect 2341 3016 2482 3019
rect 12648 3018 12653 3052
rect 12648 3017 12687 3018
rect 2356 3007 2482 3016
rect 2356 2991 2395 3007
rect 2425 2991 2482 3007
rect 2217 2969 2222 2991
rect 2284 2969 2286 2991
rect 2231 2967 2265 2969
rect 2325 2963 2434 2991
rect 2452 2969 2482 2991
rect 2515 2969 2536 2997
rect 1583 2933 1623 2959
rect 1626 2933 1643 2959
rect 1667 2955 1698 2959
rect 1725 2955 1831 2959
rect 1667 2933 1697 2955
rect 1721 2939 1831 2955
rect 1865 2945 1899 2959
rect 1947 2939 1962 2959
rect 1721 2933 1797 2939
rect 2095 2935 2125 2959
rect 2169 2935 2182 2963
rect 2452 2959 2467 2969
rect 1725 2931 1797 2933
rect 2069 2933 2135 2935
rect 2187 2933 2192 2959
rect 2314 2933 2316 2959
rect 2398 2957 2425 2959
rect 2069 2929 2101 2933
rect 2103 2929 2135 2933
rect 2324 2929 2358 2957
rect 2392 2929 2434 2957
rect 2491 2933 2536 2969
rect 2515 2929 2536 2933
rect 2549 2929 2570 3012
rect 2587 2967 2640 2990
rect 2580 2959 2640 2967
rect 2670 2987 2761 2990
rect 2670 2959 2780 2987
rect 2634 2934 2726 2936
rect 2634 2933 2681 2934
rect 1208 2911 1337 2929
rect 1443 2915 1517 2929
rect 1237 2907 1271 2911
rect 1439 2899 1517 2915
rect 1583 2923 1657 2929
rect 1583 2918 1667 2923
rect 1583 2899 1657 2918
rect 1439 2895 1491 2899
rect 1691 2897 1797 2929
rect 1846 2919 1862 2923
rect 1881 2919 1915 2929
rect 1831 2895 1947 2919
rect 1968 2918 1989 2923
rect 2043 2918 2095 2923
rect 2101 2901 2103 2929
rect 2169 2901 2216 2929
rect 2634 2925 2640 2933
rect 2670 2925 2681 2933
rect 2720 2922 2726 2934
rect 1439 2868 1457 2881
rect 1831 2868 1947 2885
rect 1208 2864 2956 2868
rect 1439 2861 1457 2864
rect 1831 2861 1947 2864
rect 1180 2836 2928 2840
rect 1142 2744 2052 2766
rect 1868 2738 1980 2744
rect 1142 2716 2052 2738
rect 1200 2652 1678 2660
rect 1868 2658 1980 2716
rect 1750 2656 2152 2658
rect 1750 2652 2120 2656
rect 230 2618 232 2628
rect 1228 2624 1678 2632
rect 1868 2630 1980 2652
rect 1750 2624 2124 2630
rect 202 2590 232 2600
rect 1868 2466 1980 2624
rect 2089 2595 2131 2607
rect 2055 2561 2161 2573
rect 2171 2509 2175 2535
rect 2255 2509 2283 2535
rect 2181 2497 2215 2509
rect 2309 2507 2325 2509
rect 2181 2475 2223 2497
rect 1879 2465 1980 2466
rect 2189 2463 2223 2475
rect 2225 2463 2233 2507
rect 2309 2463 2337 2507
rect 2349 2493 2361 2509
rect 2349 2475 2391 2493
rect 2361 2467 2391 2475
rect 2399 2489 2433 2493
rect 2445 2489 2475 2493
rect 2399 2475 2475 2489
rect 2399 2471 2433 2475
rect 2445 2467 2475 2475
rect 2115 2363 2131 2459
rect 2141 2456 2145 2457
rect 2149 2456 2165 2459
rect 2309 2457 2325 2463
rect 2361 2457 2381 2467
rect 2225 2456 2253 2457
rect 2309 2456 2339 2457
rect 2393 2456 2423 2467
rect 2445 2457 2465 2467
rect 2134 2425 2189 2456
rect 2218 2425 2293 2456
rect 2302 2425 2522 2456
rect 2134 2409 2522 2425
rect 2141 2363 2145 2409
rect 2149 2363 2165 2409
rect 2175 2395 2253 2409
rect 2265 2399 2522 2409
rect 2265 2395 2609 2399
rect 2175 2391 2609 2395
rect 2826 2393 3004 2714
rect 3682 2408 3828 2768
rect 3682 2407 3821 2408
rect 3682 2393 3708 2407
rect 2175 2383 2675 2391
rect 2175 2375 2461 2383
rect 2478 2382 2675 2383
rect 2478 2375 2491 2382
rect 2175 2363 2253 2375
rect 2283 2363 2461 2375
rect 2002 2326 2044 2344
rect 2063 2326 2501 2363
rect 2512 2348 2575 2365
rect 2632 2348 2675 2357
rect 2512 2341 2525 2348
rect 1892 2276 1912 2302
rect 1926 2276 1946 2310
rect 2002 2273 2501 2326
rect 2044 2271 2149 2272
rect 2171 2261 2391 2273
rect 2444 2261 2475 2273
rect 2171 2243 2231 2261
rect 2015 2189 2018 2243
rect 2089 2207 2141 2243
rect 2145 2211 2231 2243
rect 2233 2253 2305 2261
rect 2233 2243 2283 2253
rect 2291 2243 2299 2253
rect 2233 2211 2309 2243
rect 2325 2236 2333 2261
rect 2339 2236 2391 2261
rect 2314 2225 2406 2236
rect 2445 2225 2475 2261
rect 4438 2248 7648 2282
rect 2314 2218 2475 2225
rect 2330 2216 2475 2218
rect 2333 2211 2475 2216
rect 2145 2207 2225 2211
rect 2253 2208 2309 2211
rect 2335 2208 2475 2211
rect 2253 2207 2475 2208
rect 2095 2189 2145 2207
rect 2069 2128 2072 2189
rect 2115 2181 2145 2189
rect 2115 2177 2141 2181
rect 2149 2177 2165 2207
rect 2203 2189 2253 2207
rect 2210 2181 2253 2189
rect 2126 2174 2141 2177
rect 2210 2174 2225 2181
rect 2257 2177 2265 2207
rect 2286 2190 2434 2207
rect 2299 2189 2433 2190
rect 2294 2177 2433 2189
rect 2445 2181 2465 2207
rect 2294 2174 2309 2177
rect 2320 2171 2335 2177
rect 2320 2166 2354 2171
rect 2391 2166 2438 2171
rect 2199 2143 2377 2155
rect 2052 2112 2148 2114
rect 2199 2109 2259 2121
rect 2293 2109 2343 2121
rect 2024 2084 2120 2086
rect 1636 1972 1678 1990
rect 1750 1972 2696 1990
rect 2040 1968 2696 1972
rect 2040 1964 2592 1968
rect 1608 1944 1678 1962
rect 1750 1944 2696 1962
rect 2012 1940 2696 1944
rect 2012 1936 2620 1940
rect 1198 1866 1469 1870
rect 1534 1866 2610 1870
rect 2526 1842 2552 1848
rect 1170 1838 1469 1842
rect 1482 1834 1522 1842
rect 1534 1838 2582 1842
rect 1444 1799 1449 1811
rect 1482 1800 1541 1834
rect 403 1795 437 1799
rect -38 1614 20 1782
rect 374 1777 477 1795
rect 495 1777 529 1799
rect 543 1777 586 1795
rect 1267 1777 1365 1797
rect 1415 1777 1449 1799
rect 1507 1777 1541 1800
rect 1573 1777 1652 1805
rect 1656 1801 1658 1815
rect 1959 1801 1962 1815
rect 2526 1811 2552 1838
rect 2560 1811 2586 1814
rect 2636 1811 2666 1814
rect 2670 1811 2700 1845
rect 2740 1821 2747 1845
rect 1656 1797 1728 1801
rect 1750 1797 1836 1801
rect 1656 1783 1847 1797
rect 1849 1783 1962 1801
rect 2096 1795 2138 1801
rect 2086 1793 2138 1795
rect 1989 1783 2056 1793
rect 2085 1783 2138 1793
rect 1428 1773 1443 1777
rect 1232 1772 1262 1773
rect 340 1743 477 1761
rect 397 1739 431 1743
rect 489 1739 523 1761
rect 543 1727 552 1761
rect 562 1746 645 1772
rect 710 1746 1389 1772
rect 1417 1769 1443 1773
rect 1401 1747 1443 1769
rect 1233 1745 1365 1746
rect 1401 1745 1445 1747
rect 1238 1744 1365 1745
rect 1375 1744 1391 1745
rect 417 1719 447 1723
rect 409 1697 447 1719
rect 477 1697 527 1711
rect 409 1693 443 1697
rect 375 1659 403 1685
rect 453 1677 527 1697
rect 577 1693 586 1743
rect 590 1718 645 1744
rect 710 1733 1391 1744
rect 1401 1733 1439 1745
rect 710 1727 1439 1733
rect 620 1679 653 1713
rect 658 1680 698 1722
rect 710 1718 1403 1727
rect 1262 1713 1307 1718
rect 1320 1713 1340 1718
rect 1377 1713 1403 1718
rect 1435 1713 1439 1727
rect 1469 1713 1473 1777
rect 1520 1727 1534 1777
rect 1656 1773 1658 1783
rect 1686 1777 1762 1783
rect 1783 1777 1847 1783
rect 1848 1773 1849 1783
rect 1607 1747 1652 1771
rect 1698 1747 1700 1773
rect 1720 1747 1762 1763
rect 1812 1761 1813 1763
rect 1779 1747 1813 1761
rect 1890 1747 1891 1773
rect 1959 1747 1962 1783
rect 2185 1777 2297 1805
rect 2337 1783 2352 1801
rect 2358 1795 2424 1801
rect 2442 1799 2472 1801
rect 2427 1795 2472 1799
rect 2478 1795 2522 1801
rect 2358 1783 2522 1795
rect 2636 1783 2713 1811
rect 2358 1777 2518 1783
rect 2636 1777 2671 1783
rect 1607 1743 1813 1747
rect 1554 1727 1568 1743
rect 1644 1735 1813 1743
rect 1644 1732 1673 1735
rect 711 1679 736 1713
rect 1238 1703 1320 1713
rect 914 1699 926 1703
rect 937 1699 995 1703
rect 752 1685 804 1697
rect 834 1693 878 1697
rect 749 1679 828 1685
rect 417 1659 443 1669
rect 409 1643 443 1659
rect 453 1651 511 1677
rect 590 1666 651 1675
rect 749 1666 804 1679
rect 834 1666 889 1693
rect 914 1677 995 1699
rect 1020 1691 1142 1703
rect 1165 1695 1320 1703
rect 1363 1707 1403 1713
rect 1165 1691 1241 1695
rect 1020 1679 1241 1691
rect 409 1627 447 1643
rect 453 1627 483 1651
rect 590 1648 910 1666
rect 914 1663 1010 1677
rect 1020 1666 1142 1679
rect 1165 1668 1241 1679
rect 1262 1668 1314 1695
rect 1363 1689 1391 1707
rect 1447 1689 1473 1713
rect 1377 1679 1391 1689
rect 1454 1679 1473 1685
rect 1492 1680 1620 1727
rect 1644 1703 1658 1732
rect 1720 1727 1813 1735
rect 1644 1681 1698 1703
rect 1720 1701 1801 1727
rect 1812 1713 1813 1727
rect 1836 1732 1864 1747
rect 1915 1743 1916 1747
rect 1836 1713 1849 1732
rect 1815 1703 1849 1713
rect 1881 1709 1916 1713
rect 1922 1709 1977 1747
rect 1985 1743 2041 1747
rect 2086 1743 2120 1747
rect 2033 1724 2085 1739
rect 1959 1703 1977 1709
rect 1815 1701 1890 1703
rect 1914 1701 1977 1703
rect 1980 1713 2014 1717
rect 2033 1713 2050 1724
rect 1980 1709 2050 1713
rect 1728 1691 1774 1701
rect 1741 1689 1774 1691
rect 1815 1689 1978 1701
rect 1744 1681 1774 1689
rect 1165 1666 1314 1668
rect 1320 1666 1340 1679
rect 1354 1666 1366 1679
rect 1377 1666 1400 1679
rect 1439 1666 1454 1679
rect 1473 1675 1488 1679
rect 1459 1666 1488 1675
rect 1513 1666 1528 1680
rect 1539 1675 1620 1680
rect 1641 1675 1698 1681
rect 1728 1679 1774 1681
rect 1830 1679 1978 1689
rect 1744 1678 1774 1679
rect 1539 1666 1698 1675
rect 1020 1663 1698 1666
rect 1729 1663 1789 1678
rect 1812 1663 1813 1679
rect 1830 1667 1890 1679
rect 1914 1675 1978 1679
rect 1980 1675 2014 1709
rect 2033 1675 2050 1709
rect 2056 1675 2085 1724
rect 2185 1713 2188 1777
rect 2201 1773 2216 1777
rect 2201 1771 2227 1773
rect 2283 1771 2304 1773
rect 2201 1747 2304 1771
rect 2358 1747 2364 1777
rect 2382 1751 2388 1773
rect 2492 1772 2518 1777
rect 2449 1761 2582 1772
rect 2392 1747 2582 1761
rect 2219 1743 2298 1747
rect 2219 1713 2222 1743
rect 2253 1737 2298 1743
rect 2253 1713 2254 1737
rect 2337 1732 2364 1747
rect 2387 1746 2582 1747
rect 2703 1746 2713 1783
rect 2387 1744 2534 1746
rect 2387 1735 2610 1744
rect 2352 1713 2364 1732
rect 2392 1713 2398 1735
rect 2403 1727 2610 1735
rect 2424 1718 2610 1727
rect 2424 1713 2518 1718
rect 2522 1717 2534 1718
rect 2086 1709 2120 1713
rect 2253 1703 2298 1713
rect 2253 1699 2254 1703
rect 2253 1691 2274 1699
rect 2086 1675 2132 1691
rect 2201 1684 2219 1691
rect 2253 1684 2291 1691
rect 1914 1667 1977 1675
rect 1830 1663 1978 1667
rect 989 1649 1010 1663
rect 591 1647 611 1648
rect 409 1625 483 1627
rect 443 1609 483 1625
rect 565 1638 623 1647
rect 749 1638 759 1648
rect 783 1645 828 1648
rect 783 1643 793 1645
rect 804 1643 825 1645
rect 783 1638 835 1643
rect 862 1642 895 1648
rect 565 1624 910 1638
rect 968 1631 977 1649
rect 980 1634 1020 1649
rect 989 1631 1020 1634
rect 562 1620 910 1624
rect 453 1598 483 1609
rect 447 1593 483 1598
rect -17 1559 114 1587
rect 147 1571 369 1583
rect 443 1575 483 1593
rect 207 1559 369 1571
rect 447 1568 483 1575
rect 522 1570 523 1613
rect 577 1607 611 1620
rect 749 1607 759 1620
rect 783 1607 793 1620
rect 669 1595 793 1607
rect 804 1617 861 1620
rect 447 1559 450 1568
rect 512 1561 523 1570
rect 539 1569 565 1593
rect 623 1569 649 1593
rect 668 1576 796 1595
rect 804 1593 834 1617
rect 955 1607 1020 1631
rect 804 1583 861 1593
rect 804 1581 834 1583
rect 804 1576 841 1581
rect 461 1559 523 1561
rect 668 1561 841 1576
rect 880 1571 946 1597
rect 968 1587 977 1607
rect 989 1593 1020 1607
rect 1023 1593 1044 1663
rect 1110 1659 1655 1663
rect 1698 1659 1717 1663
rect 1744 1659 1770 1663
rect 1060 1645 1091 1657
rect 1110 1652 1770 1659
rect 1806 1652 1816 1663
rect 1846 1652 1847 1663
rect 1881 1652 1986 1663
rect 1110 1650 2002 1652
rect 2007 1650 2085 1675
rect 2115 1657 2136 1675
rect 2086 1650 2136 1657
rect 2177 1668 2182 1684
rect 2201 1679 2291 1684
rect 2201 1675 2274 1679
rect 2185 1668 2201 1675
rect 2212 1668 2274 1675
rect 2333 1669 2336 1691
rect 2352 1669 2358 1713
rect 2367 1689 2401 1713
rect 2424 1701 2515 1713
rect 2424 1685 2492 1701
rect 2437 1679 2492 1685
rect 2177 1657 2274 1668
rect 2302 1657 2333 1669
rect 2336 1659 2367 1669
rect 2398 1659 2428 1675
rect 2437 1659 2458 1679
rect 2522 1675 2552 1717
rect 2630 1685 2646 1717
rect 2702 1696 2713 1746
rect 3682 1752 3844 2224
rect 6107 2180 6108 2234
rect 6161 2159 6162 2180
rect 6173 2159 7549 2168
rect 6074 2125 6085 2136
rect 6097 2125 6108 2136
rect 6157 2134 7565 2159
rect 7606 2136 7615 2234
rect 6161 2128 6246 2134
rect 7457 2128 7561 2134
rect 6161 2125 6210 2128
rect 7457 2126 7538 2128
rect 7457 2125 7552 2126
rect 7606 2125 7617 2136
rect 7629 2125 7640 2136
rect 6074 2059 6108 2125
rect 6160 2122 6226 2125
rect 7457 2122 7554 2125
rect 6133 2100 6218 2122
rect 7457 2109 7552 2122
rect 7606 2121 7640 2125
rect 7496 2100 7552 2109
rect 7602 2109 7648 2121
rect 6176 2084 6210 2100
rect 7504 2084 7538 2100
rect 6074 2048 6085 2059
rect 6097 2048 6108 2059
rect 6133 2062 6218 2084
rect 7496 2062 7552 2084
rect 7602 2075 7640 2109
rect 7602 2063 7648 2075
rect 6133 1982 6144 2062
rect 6160 2059 6226 2062
rect 7488 2059 7554 2062
rect 7606 2059 7640 2063
rect 6161 2056 6176 2059
rect 7496 2058 7552 2059
rect 6161 2050 6246 2056
rect 7468 2050 7561 2056
rect 6157 2025 7565 2050
rect 7606 2048 7617 2059
rect 7629 2048 7640 2059
rect 6161 2010 6172 2025
rect 6173 2016 7549 2025
rect 6161 2004 6162 2010
rect 7606 2004 7615 2048
rect 8902 1978 9106 1980
rect 4438 1902 7648 1936
rect 3682 1728 3862 1752
rect 8196 1750 8224 1752
rect 3682 1724 3844 1728
rect 3682 1700 3890 1724
rect 2679 1685 2690 1686
rect 2585 1679 2690 1685
rect 2490 1667 2520 1675
rect 2522 1667 2534 1675
rect 2471 1659 2534 1667
rect 2336 1657 2534 1659
rect 2177 1654 2291 1657
rect 2177 1650 2232 1654
rect 2253 1650 2291 1654
rect 2304 1650 2331 1657
rect 2333 1650 2336 1657
rect 2352 1656 2358 1657
rect 2363 1656 2534 1657
rect 2348 1650 2534 1656
rect 1110 1649 2534 1650
rect 2574 1654 2594 1675
rect 2630 1654 2646 1679
rect 2679 1675 2690 1679
rect 2702 1685 2721 1696
rect 2679 1671 2688 1675
rect 2702 1671 2713 1685
rect 2679 1654 2713 1671
rect 2574 1649 2713 1654
rect 2727 1649 2742 1663
rect 1110 1648 2567 1649
rect 2579 1648 2750 1649
rect 1125 1645 1366 1648
rect 1142 1638 1180 1645
rect 1183 1638 1366 1645
rect 1377 1638 1400 1648
rect 1454 1645 1473 1648
rect 1513 1638 1530 1648
rect 1547 1647 1573 1648
rect 1581 1647 1744 1648
rect 1547 1641 1745 1647
rect 1774 1645 1830 1648
rect 1846 1646 1847 1648
rect 1875 1646 2028 1648
rect 1567 1638 1745 1641
rect 1110 1634 1745 1638
rect 1110 1631 1694 1634
rect 1698 1631 1745 1634
rect 1110 1629 1745 1631
rect 1098 1627 1745 1629
rect 1094 1624 1745 1627
rect 1770 1624 1830 1645
rect 1841 1641 2028 1646
rect 1841 1637 2018 1641
rect 1841 1634 2012 1637
rect 1841 1627 1969 1634
rect 1841 1624 1972 1627
rect 1973 1624 2003 1634
rect 2041 1625 2085 1648
rect 2086 1641 2132 1648
rect 2177 1637 2232 1648
rect 2253 1645 2291 1648
rect 2304 1641 2331 1648
rect 1094 1623 2003 1624
rect 1098 1622 2003 1623
rect 2056 1622 2094 1625
rect 2141 1623 2232 1637
rect 2274 1623 2301 1639
rect 2333 1635 2336 1648
rect 2348 1637 2567 1648
rect 2141 1622 2253 1623
rect 2257 1622 2301 1623
rect 2348 1633 2520 1637
rect 2522 1634 2564 1637
rect 2615 1634 2750 1648
rect 2802 1635 2830 1699
rect 3204 1677 3248 1699
rect 2836 1635 2864 1665
rect 2522 1633 2560 1634
rect 2348 1630 2580 1633
rect 2348 1629 2604 1630
rect 2348 1627 2614 1629
rect 2630 1627 2716 1634
rect 2348 1626 2620 1627
rect 2625 1626 2716 1627
rect 2348 1622 2716 1626
rect 1098 1620 2716 1622
rect 991 1587 1025 1593
rect 965 1583 1025 1587
rect 1048 1583 1050 1597
rect 1098 1593 1366 1620
rect 1377 1593 1400 1620
rect 1429 1617 1448 1620
rect 1454 1617 1481 1620
rect 1429 1593 1454 1617
rect 1481 1593 1488 1617
rect 1094 1591 1354 1593
rect 1094 1590 1351 1591
rect 1094 1589 1340 1590
rect 1142 1585 1311 1589
rect 1142 1583 1301 1585
rect 917 1569 933 1571
rect 965 1565 1036 1583
rect 1048 1579 1120 1583
rect 1142 1579 1351 1583
rect 1359 1580 1392 1593
rect 1454 1583 1481 1593
rect 1528 1589 1530 1620
rect 1579 1619 1830 1620
rect 1579 1614 1779 1619
rect 1806 1614 1830 1619
rect 1841 1614 1972 1620
rect 1579 1607 1972 1614
rect 1973 1607 2003 1620
rect 2056 1613 2136 1620
rect 2141 1613 2253 1620
rect 1532 1593 1558 1597
rect 1600 1593 1969 1607
rect 1972 1604 2003 1607
rect 2006 1604 2028 1607
rect 2056 1604 2253 1613
rect 2257 1608 2301 1620
rect 2348 1609 2620 1620
rect 2358 1608 2620 1609
rect 2257 1604 2620 1608
rect 1972 1594 2620 1604
rect 1972 1593 2003 1594
rect 1532 1589 1577 1593
rect 1528 1583 1577 1589
rect 1359 1579 1406 1580
rect 1414 1579 1429 1580
rect 1048 1576 1354 1579
rect 1048 1565 1239 1576
rect 1241 1565 1354 1576
rect 668 1560 861 1561
rect 705 1559 861 1560
rect 965 1559 1023 1565
rect 17 1525 80 1553
rect 288 1549 309 1555
rect 207 1536 335 1549
rect 387 1548 417 1555
rect 443 1548 523 1559
rect 342 1539 523 1548
rect 530 1539 542 1559
rect 564 1539 576 1559
rect 342 1536 576 1539
rect 207 1530 576 1536
rect 624 1530 654 1555
rect 705 1545 753 1559
rect 757 1545 835 1559
rect 705 1539 835 1545
rect 861 1539 865 1559
rect 912 1539 926 1559
rect 705 1530 937 1539
rect -17 1427 3 1525
rect 17 1427 37 1525
rect 144 1514 162 1529
rect 207 1528 937 1530
rect 955 1529 960 1559
rect 965 1529 989 1559
rect 1048 1555 1050 1565
rect 1078 1559 1154 1565
rect 1129 1555 1154 1559
rect 1156 1555 1239 1565
rect 1240 1555 1307 1565
rect 999 1529 1023 1553
rect 1090 1529 1092 1555
rect 1112 1539 1154 1545
rect 1182 1543 1232 1555
rect 1282 1546 1312 1555
rect 1171 1539 1232 1543
rect 1112 1531 1221 1539
rect 1112 1530 1239 1531
rect 1273 1530 1307 1531
rect 1351 1530 1354 1565
rect 1359 1565 1448 1579
rect 1488 1577 1577 1583
rect 1478 1575 1577 1577
rect 1477 1569 1577 1575
rect 1600 1580 1972 1593
rect 1973 1580 2003 1593
rect 2006 1587 2028 1594
rect 2056 1593 2620 1594
rect 2056 1589 2380 1593
rect 1600 1576 2018 1580
rect 2052 1576 2380 1589
rect 2388 1591 2620 1593
rect 2388 1576 2458 1591
rect 2471 1576 2620 1591
rect 1600 1573 2620 1576
rect 1600 1570 1675 1573
rect 1477 1565 1558 1569
rect 1359 1559 1392 1565
rect 1406 1549 1425 1565
rect 1429 1564 1433 1565
rect 1528 1555 1558 1565
rect 1593 1565 1675 1570
rect 1593 1559 1608 1565
rect 1616 1559 1675 1565
rect 1688 1565 2620 1573
rect 1688 1559 1774 1565
rect 1784 1559 1912 1565
rect 1921 1559 2062 1565
rect 1391 1534 1448 1549
rect 1528 1539 1549 1555
rect 1573 1553 1645 1559
rect 1688 1555 1729 1559
rect 1675 1553 1729 1555
rect 1573 1539 1729 1553
rect 1406 1530 1425 1534
rect 1528 1530 1729 1539
rect 1110 1529 1729 1530
rect 1744 1555 1774 1559
rect 1779 1555 1822 1559
rect 1744 1551 1822 1555
rect 1744 1533 1834 1551
rect 1878 1549 1912 1559
rect 1744 1529 1829 1533
rect 1850 1531 1876 1543
rect 1884 1531 1912 1549
rect 1850 1529 1884 1531
rect 1897 1529 1912 1531
rect 1925 1557 2062 1559
rect 2101 1559 2620 1565
rect 2625 1577 2716 1620
rect 2625 1561 2674 1577
rect 2101 1557 2472 1559
rect 1925 1529 2085 1557
rect 207 1525 335 1528
rect 226 1514 246 1525
rect 319 1515 339 1525
rect 144 1499 147 1514
rect 136 1496 186 1499
rect 226 1496 231 1514
rect 267 1496 270 1515
rect 301 1508 304 1515
rect 329 1508 339 1515
rect 359 1508 542 1528
rect 286 1502 542 1508
rect 557 1514 582 1528
rect 625 1527 654 1528
rect 669 1515 696 1527
rect 705 1526 937 1528
rect 705 1525 757 1526
rect 705 1515 753 1525
rect 767 1517 937 1526
rect 950 1525 1023 1529
rect 1036 1527 1675 1529
rect 1696 1527 1756 1529
rect 1779 1527 2085 1529
rect 2101 1547 2380 1557
rect 2388 1547 2415 1557
rect 2442 1547 2470 1557
rect 2481 1549 2620 1559
rect 2481 1547 2583 1549
rect 2101 1527 2398 1547
rect 2442 1527 2472 1547
rect 2481 1527 2490 1547
rect 2520 1543 2583 1547
rect 2596 1543 2617 1549
rect 2520 1533 2574 1543
rect 2630 1527 2674 1561
rect 2679 1569 2708 1577
rect 2721 1569 2750 1634
rect 3049 1631 3083 1665
rect 3170 1643 3248 1665
rect 3282 1631 3296 1665
rect 3316 1659 3330 1699
rect 3682 1674 3844 1700
rect 3682 1673 3825 1674
rect 3682 1672 3712 1673
rect 3682 1631 3698 1672
rect 2761 1569 2776 1629
rect 2915 1601 2928 1629
rect 2873 1597 3009 1601
rect 2873 1589 3015 1597
rect 2873 1585 2928 1589
rect 2828 1569 2830 1585
rect 2862 1569 2864 1585
rect 2873 1569 2925 1585
rect 2949 1573 3015 1589
rect 3030 1573 3097 1628
rect 3183 1601 3214 1631
rect 3217 1615 3248 1631
rect 3217 1601 3334 1615
rect 3123 1597 3143 1601
rect 3155 1600 3177 1601
rect 3180 1600 3334 1601
rect 3117 1586 3143 1597
rect 3117 1573 3131 1586
rect 3146 1580 3334 1600
rect 3146 1573 3177 1580
rect 3183 1573 3334 1580
rect 2679 1554 2888 1569
rect 2679 1527 2873 1554
rect 2909 1527 2925 1569
rect 2928 1527 3334 1573
rect 557 1502 576 1514
rect 623 1502 630 1511
rect 657 1502 664 1511
rect 669 1510 699 1515
rect 705 1510 706 1515
rect 669 1502 706 1510
rect 769 1512 937 1517
rect 769 1503 839 1512
rect 851 1511 865 1512
rect 887 1511 937 1512
rect 851 1509 937 1511
rect 946 1509 1006 1525
rect 1036 1517 3334 1527
rect 1036 1514 1065 1517
rect 769 1502 783 1503
rect 792 1502 831 1503
rect 851 1502 1012 1509
rect 286 1500 1012 1502
rect 301 1496 304 1500
rect 329 1497 339 1500
rect 359 1499 542 1500
rect 318 1496 339 1497
rect 136 1467 359 1496
rect 144 1465 157 1467
rect 102 1460 157 1465
rect 170 1465 359 1467
rect 406 1480 542 1499
rect 406 1470 527 1480
rect 406 1465 496 1470
rect 170 1461 387 1465
rect 417 1461 462 1465
rect 170 1460 462 1461
rect 102 1445 162 1460
rect 170 1450 465 1460
rect 170 1449 387 1450
rect 201 1445 298 1449
rect 301 1445 304 1449
rect 318 1445 387 1449
rect 392 1449 415 1450
rect 417 1449 465 1450
rect 483 1449 496 1465
rect 392 1445 527 1449
rect 102 1433 155 1445
rect 189 1433 387 1445
rect 141 1427 155 1433
rect 175 1429 387 1433
rect 393 1429 527 1445
rect 530 1439 542 1480
rect 557 1473 576 1500
rect 623 1477 630 1500
rect 654 1495 706 1500
rect 557 1460 567 1473
rect 654 1470 699 1495
rect 753 1494 1012 1500
rect 1036 1494 1050 1514
rect 1110 1512 3334 1517
rect 1112 1503 3334 1512
rect 1112 1502 1193 1503
rect 1199 1502 3334 1503
rect 753 1475 1057 1494
rect 1110 1484 3334 1502
rect 1112 1483 3334 1484
rect 654 1460 666 1470
rect 769 1467 783 1475
rect 792 1467 1057 1475
rect 557 1449 582 1460
rect 654 1457 681 1460
rect 698 1457 706 1463
rect 654 1449 706 1457
rect 557 1448 612 1449
rect 619 1448 708 1449
rect 557 1445 708 1448
rect 175 1427 527 1429
rect -17 1422 527 1427
rect -17 1407 387 1422
rect 393 1411 527 1422
rect 392 1407 527 1411
rect 582 1417 612 1445
rect 619 1417 708 1445
rect 582 1407 708 1417
rect 749 1407 758 1467
rect 769 1453 1057 1467
rect 1101 1475 3334 1483
rect 1101 1467 1179 1475
rect 769 1433 827 1453
rect 851 1449 1057 1453
rect 1060 1449 1086 1457
rect 1101 1449 1120 1467
rect 1149 1460 1179 1467
rect 1182 1460 3334 1475
rect 1134 1453 3334 1460
rect 1134 1449 1194 1453
rect 1199 1449 3334 1453
rect 851 1445 1090 1449
rect 851 1437 905 1445
rect 920 1437 960 1445
rect 976 1437 999 1445
rect 1026 1437 1033 1445
rect 1046 1437 1090 1445
rect 769 1407 821 1433
rect 849 1407 1090 1437
rect 1101 1429 3334 1449
rect 8902 1434 8907 1468
rect 8902 1433 8941 1434
rect 1111 1413 3334 1429
rect 1111 1407 2523 1413
rect -17 1387 2523 1407
rect 2577 1395 2606 1413
rect 2721 1398 2730 1413
rect 2584 1387 2606 1395
rect 2618 1392 2710 1398
rect 2618 1387 2699 1392
rect 2798 1391 3334 1413
rect -17 1381 2520 1387
rect -7 1359 2520 1381
rect 35 1353 2520 1359
rect 35 1351 2523 1353
rect 2584 1351 2606 1353
rect 35 1326 2526 1351
rect 2618 1329 2688 1387
rect 2710 1353 2776 1372
rect 2798 1365 2818 1391
rect 2828 1369 2949 1387
rect 2996 1369 3138 1387
rect 3172 1369 3217 1387
rect 2710 1329 2742 1338
rect -272 1293 -233 1325
rect 35 1324 2610 1326
rect 2618 1324 2742 1329
rect 35 1322 2742 1324
rect 35 1298 2526 1322
rect 2618 1319 2742 1322
rect 2530 1298 2560 1317
rect 35 1296 2582 1298
rect 2598 1296 2614 1301
rect 2618 1296 2710 1319
rect 35 1294 2728 1296
rect 35 1293 2526 1294
rect 97 1292 117 1293
rect 147 1292 201 1293
rect 184 1290 201 1292
rect -28 1256 38 1276
rect 169 1275 201 1290
rect 214 1284 238 1293
rect 243 1284 266 1293
rect 184 1249 189 1275
rect 214 1256 231 1284
rect 279 1281 313 1293
rect 333 1281 417 1293
rect 279 1276 347 1281
rect 238 1256 243 1276
rect 279 1273 374 1276
rect 257 1267 374 1273
rect 443 1269 452 1293
rect 453 1271 483 1293
rect 418 1267 443 1269
rect 452 1267 477 1269
rect 257 1259 440 1267
rect 443 1259 452 1267
rect 522 1259 523 1293
rect 543 1285 645 1293
rect 543 1269 608 1285
rect 659 1283 696 1293
rect 709 1283 741 1293
rect 749 1283 758 1293
rect 787 1283 822 1293
rect 825 1283 827 1293
rect 617 1273 683 1283
rect 699 1279 835 1283
rect 257 1256 452 1259
rect 543 1257 608 1267
rect 617 1257 695 1273
rect 699 1268 753 1279
rect 783 1271 835 1279
rect 783 1268 792 1271
rect 822 1268 835 1271
rect 214 1251 238 1256
rect 215 1248 238 1251
rect 243 1248 452 1256
rect 0 1228 38 1248
rect 238 1228 243 1248
rect 257 1247 452 1248
rect 299 1239 374 1247
rect 381 1239 452 1247
rect 299 1235 452 1239
rect 300 1233 452 1235
rect 495 1233 529 1257
rect 543 1235 695 1257
rect 587 1233 695 1235
rect 709 1267 753 1268
rect 787 1267 792 1268
rect 825 1267 827 1268
rect 859 1267 861 1293
rect 901 1283 1033 1293
rect 901 1281 1035 1283
rect 887 1271 1035 1281
rect 903 1268 932 1271
rect 941 1269 1035 1271
rect 903 1267 918 1268
rect 709 1245 792 1267
rect 901 1261 935 1267
rect 709 1233 753 1245
rect 300 1229 381 1233
rect 300 1228 418 1229
rect 300 1217 313 1228
rect 352 1221 418 1228
rect 381 1217 418 1221
rect 617 1219 719 1233
rect 217 1215 247 1217
rect 381 1199 452 1217
rect 397 1195 431 1199
rect 489 1183 523 1217
rect 527 1203 561 1219
rect 599 1203 719 1219
rect 527 1199 719 1203
rect 527 1185 721 1199
rect 669 1173 685 1185
rect 693 1173 721 1185
rect 693 1169 719 1173
rect 735 1169 759 1233
rect 787 1199 793 1233
rect 825 1221 827 1233
rect 829 1199 835 1261
rect 901 1241 939 1261
rect 859 1203 861 1233
rect 867 1203 873 1223
rect 903 1214 939 1241
rect 953 1237 1035 1269
rect 1039 1267 1067 1293
rect 1149 1289 1179 1293
rect 1198 1289 1221 1293
rect 1069 1271 1088 1283
rect 1149 1271 1175 1289
rect 1193 1282 1221 1289
rect 1289 1283 1293 1293
rect 1311 1283 2526 1293
rect 1187 1271 1221 1282
rect 1247 1280 2526 1283
rect 1247 1273 1569 1280
rect 1229 1271 1569 1273
rect 1069 1268 1334 1271
rect 1338 1268 1353 1271
rect 1421 1268 1437 1271
rect 1069 1256 1275 1268
rect 1069 1245 1179 1256
rect 1187 1248 1275 1256
rect 953 1221 1007 1237
rect 1090 1233 1103 1245
rect 1073 1225 1103 1233
rect 953 1217 983 1221
rect 1049 1217 1103 1225
rect 1107 1239 1179 1245
rect 1193 1239 1199 1248
rect 1203 1239 1275 1248
rect 1107 1233 1265 1239
rect 1107 1219 1247 1233
rect 1289 1228 1319 1268
rect 1436 1243 1437 1268
rect 1446 1247 1569 1271
rect 1593 1267 1598 1280
rect 1599 1271 1665 1280
rect 1599 1267 1668 1271
rect 1699 1267 1715 1280
rect 1738 1271 1740 1280
rect 1723 1267 1782 1271
rect 1807 1267 1884 1280
rect 1903 1271 1942 1280
rect 1927 1268 1942 1271
rect 1974 1267 2526 1280
rect 2530 1267 2560 1294
rect 2598 1283 2614 1294
rect 1467 1243 1569 1247
rect 1399 1233 1569 1243
rect 1599 1259 1699 1267
rect 1329 1228 1344 1233
rect 1436 1231 1437 1233
rect 1467 1231 1569 1233
rect 1477 1228 1507 1231
rect 1559 1228 1564 1231
rect 1593 1228 1598 1233
rect 1599 1231 1668 1259
rect 1723 1256 1864 1267
rect 1897 1257 2510 1267
rect 2564 1258 2582 1267
rect 2598 1258 2616 1283
rect 1738 1247 1864 1256
rect 1738 1231 1777 1247
rect 1807 1231 1864 1247
rect 1599 1228 1604 1231
rect 1666 1228 1668 1231
rect 1707 1228 1816 1231
rect 1834 1228 1864 1231
rect 1897 1233 1952 1252
rect 1974 1245 2510 1257
rect 2011 1233 2195 1245
rect 1897 1228 1918 1233
rect 1931 1228 1952 1233
rect 2049 1228 2121 1233
rect 2141 1228 2195 1233
rect 2249 1233 2383 1245
rect 2249 1228 2301 1233
rect 2309 1228 2388 1233
rect 2393 1228 2422 1233
rect 2618 1228 2710 1294
rect 1107 1217 1281 1219
rect 1289 1217 2924 1228
rect 953 1214 2924 1217
rect 903 1206 2924 1214
rect 769 1169 793 1199
rect 859 1173 899 1203
rect 903 1202 2582 1206
rect 903 1200 1522 1202
rect 1551 1200 1564 1202
rect 1834 1200 1849 1202
rect 1873 1200 1918 1202
rect 1931 1200 1952 1202
rect 1995 1200 2489 1202
rect 903 1199 2896 1200
rect 965 1173 1005 1199
rect 1008 1173 1025 1199
rect 1049 1195 1080 1199
rect 1107 1195 1213 1199
rect 1049 1173 1079 1195
rect 1103 1179 1213 1195
rect 1247 1185 1281 1199
rect 1103 1173 1179 1179
rect 1293 1178 2896 1199
rect 1293 1174 2610 1178
rect 1107 1171 1179 1173
rect 1451 1173 1517 1174
rect 1569 1173 1574 1174
rect 1696 1173 1698 1174
rect 1451 1169 1483 1173
rect 1485 1169 1517 1173
rect 1706 1169 1740 1174
rect 1774 1169 1816 1174
rect 1873 1173 1918 1174
rect 1897 1169 1918 1173
rect 1931 1169 1952 1174
rect 2301 1173 2331 1174
rect 2353 1173 2388 1174
rect 2359 1169 2388 1173
rect 2393 1173 2425 1174
rect 2393 1169 2422 1173
rect 590 1151 719 1169
rect 825 1155 899 1169
rect 619 1147 653 1151
rect 821 1139 899 1155
rect 965 1163 1039 1169
rect 965 1158 1049 1163
rect 965 1139 1039 1158
rect 821 1135 873 1139
rect 1073 1137 1179 1169
rect 1228 1159 1244 1163
rect 1263 1159 1297 1169
rect 1213 1135 1329 1159
rect 1350 1158 1371 1163
rect 1425 1158 1477 1163
rect 1483 1141 1485 1169
rect 1551 1141 1598 1169
rect 1999 1165 2341 1169
rect 2049 1158 2067 1161
rect 2131 1158 2158 1161
rect 2299 1158 2346 1161
rect 2383 1158 2435 1161
rect 821 1108 839 1121
rect 1213 1108 1329 1125
rect 590 1104 2002 1108
rect 821 1101 839 1104
rect 1213 1101 1329 1104
rect 562 1076 1974 1080
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use int_pfd_cp  int_pfd_cp_0
timestamp 1708427081
transform 1 0 824 0 1 6024
box -1298 -8024 13490 10103
use int_pfd_cp  int_pfd_cp_1
timestamp 1708427081
transform 1 0 862 0 1 6024
box -1298 -8024 13490 10103
use int_pfd_cp  int_pfd_cp_2
timestamp 1708427081
transform 1 0 1298 0 1 8624
box -1298 -8024 13490 10103
use int_pfd_cp  x1
timestamp 1708427081
transform 1 0 0 0 1 600
box -1298 -8024 13490 10103
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 cp_bias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 A
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 B
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 cp_out
port 5 nsew
<< end >>
