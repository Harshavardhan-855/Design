magic
tech sky130A
magscale 1 2
timestamp 1706788245
<< error_p >>
rect -560 5072 -502 5078
rect -442 5072 -384 5078
rect -324 5072 -266 5078
rect -206 5072 -148 5078
rect -88 5072 -30 5078
rect 30 5072 88 5078
rect 148 5072 206 5078
rect 266 5072 324 5078
rect 384 5072 442 5078
rect 502 5072 560 5078
rect -560 5038 -548 5072
rect -442 5038 -430 5072
rect -324 5038 -312 5072
rect -206 5038 -194 5072
rect -88 5038 -76 5072
rect 30 5038 42 5072
rect 148 5038 160 5072
rect 266 5038 278 5072
rect 384 5038 396 5072
rect 502 5038 514 5072
rect -560 5032 -502 5038
rect -442 5032 -384 5038
rect -324 5032 -266 5038
rect -206 5032 -148 5038
rect -88 5032 -30 5038
rect 30 5032 88 5038
rect 148 5032 206 5038
rect 266 5032 324 5038
rect 384 5032 442 5038
rect 502 5032 560 5038
rect -560 -5038 -502 -5032
rect -442 -5038 -384 -5032
rect -324 -5038 -266 -5032
rect -206 -5038 -148 -5032
rect -88 -5038 -30 -5032
rect 30 -5038 88 -5032
rect 148 -5038 206 -5032
rect 266 -5038 324 -5032
rect 384 -5038 442 -5032
rect 502 -5038 560 -5032
rect -560 -5072 -548 -5038
rect -442 -5072 -430 -5038
rect -324 -5072 -312 -5038
rect -206 -5072 -194 -5038
rect -88 -5072 -76 -5038
rect 30 -5072 42 -5038
rect 148 -5072 160 -5038
rect 266 -5072 278 -5038
rect 384 -5072 396 -5038
rect 502 -5072 514 -5038
rect -560 -5078 -502 -5072
rect -442 -5078 -384 -5072
rect -324 -5078 -266 -5072
rect -206 -5078 -148 -5072
rect -88 -5078 -30 -5072
rect 30 -5078 88 -5072
rect 148 -5078 206 -5072
rect 266 -5078 324 -5072
rect 384 -5078 442 -5072
rect 502 -5078 560 -5072
<< pwell >>
rect -757 -5210 757 5210
<< nmos >>
rect -561 -5000 -501 5000
rect -443 -5000 -383 5000
rect -325 -5000 -265 5000
rect -207 -5000 -147 5000
rect -89 -5000 -29 5000
rect 29 -5000 89 5000
rect 147 -5000 207 5000
rect 265 -5000 325 5000
rect 383 -5000 443 5000
rect 501 -5000 561 5000
<< ndiff >>
rect -619 4988 -561 5000
rect -619 -4988 -607 4988
rect -573 -4988 -561 4988
rect -619 -5000 -561 -4988
rect -501 4988 -443 5000
rect -501 -4988 -489 4988
rect -455 -4988 -443 4988
rect -501 -5000 -443 -4988
rect -383 4988 -325 5000
rect -383 -4988 -371 4988
rect -337 -4988 -325 4988
rect -383 -5000 -325 -4988
rect -265 4988 -207 5000
rect -265 -4988 -253 4988
rect -219 -4988 -207 4988
rect -265 -5000 -207 -4988
rect -147 4988 -89 5000
rect -147 -4988 -135 4988
rect -101 -4988 -89 4988
rect -147 -5000 -89 -4988
rect -29 4988 29 5000
rect -29 -4988 -17 4988
rect 17 -4988 29 4988
rect -29 -5000 29 -4988
rect 89 4988 147 5000
rect 89 -4988 101 4988
rect 135 -4988 147 4988
rect 89 -5000 147 -4988
rect 207 4988 265 5000
rect 207 -4988 219 4988
rect 253 -4988 265 4988
rect 207 -5000 265 -4988
rect 325 4988 383 5000
rect 325 -4988 337 4988
rect 371 -4988 383 4988
rect 325 -5000 383 -4988
rect 443 4988 501 5000
rect 443 -4988 455 4988
rect 489 -4988 501 4988
rect 443 -5000 501 -4988
rect 561 4988 619 5000
rect 561 -4988 573 4988
rect 607 -4988 619 4988
rect 561 -5000 619 -4988
<< ndiffc >>
rect -607 -4988 -573 4988
rect -489 -4988 -455 4988
rect -371 -4988 -337 4988
rect -253 -4988 -219 4988
rect -135 -4988 -101 4988
rect -17 -4988 17 4988
rect 101 -4988 135 4988
rect 219 -4988 253 4988
rect 337 -4988 371 4988
rect 455 -4988 489 4988
rect 573 -4988 607 4988
<< psubdiff >>
rect -721 5140 -625 5174
rect 625 5140 721 5174
rect -721 5078 -687 5140
rect 687 5078 721 5140
rect -721 -5140 -687 -5078
rect 687 -5140 721 -5078
rect -721 -5174 -625 -5140
rect 625 -5174 721 -5140
<< psubdiffcont >>
rect -625 5140 625 5174
rect -721 -5078 -687 5078
rect 687 -5078 721 5078
rect -625 -5174 625 -5140
<< poly >>
rect -564 5072 -498 5088
rect -564 5038 -548 5072
rect -514 5038 -498 5072
rect -564 5022 -498 5038
rect -446 5072 -380 5088
rect -446 5038 -430 5072
rect -396 5038 -380 5072
rect -446 5022 -380 5038
rect -328 5072 -262 5088
rect -328 5038 -312 5072
rect -278 5038 -262 5072
rect -328 5022 -262 5038
rect -210 5072 -144 5088
rect -210 5038 -194 5072
rect -160 5038 -144 5072
rect -210 5022 -144 5038
rect -92 5072 -26 5088
rect -92 5038 -76 5072
rect -42 5038 -26 5072
rect -92 5022 -26 5038
rect 26 5072 92 5088
rect 26 5038 42 5072
rect 76 5038 92 5072
rect 26 5022 92 5038
rect 144 5072 210 5088
rect 144 5038 160 5072
rect 194 5038 210 5072
rect 144 5022 210 5038
rect 262 5072 328 5088
rect 262 5038 278 5072
rect 312 5038 328 5072
rect 262 5022 328 5038
rect 380 5072 446 5088
rect 380 5038 396 5072
rect 430 5038 446 5072
rect 380 5022 446 5038
rect 498 5072 564 5088
rect 498 5038 514 5072
rect 548 5038 564 5072
rect 498 5022 564 5038
rect -561 5000 -501 5022
rect -443 5000 -383 5022
rect -325 5000 -265 5022
rect -207 5000 -147 5022
rect -89 5000 -29 5022
rect 29 5000 89 5022
rect 147 5000 207 5022
rect 265 5000 325 5022
rect 383 5000 443 5022
rect 501 5000 561 5022
rect -561 -5022 -501 -5000
rect -443 -5022 -383 -5000
rect -325 -5022 -265 -5000
rect -207 -5022 -147 -5000
rect -89 -5022 -29 -5000
rect 29 -5022 89 -5000
rect 147 -5022 207 -5000
rect 265 -5022 325 -5000
rect 383 -5022 443 -5000
rect 501 -5022 561 -5000
rect -564 -5038 -498 -5022
rect -564 -5072 -548 -5038
rect -514 -5072 -498 -5038
rect -564 -5088 -498 -5072
rect -446 -5038 -380 -5022
rect -446 -5072 -430 -5038
rect -396 -5072 -380 -5038
rect -446 -5088 -380 -5072
rect -328 -5038 -262 -5022
rect -328 -5072 -312 -5038
rect -278 -5072 -262 -5038
rect -328 -5088 -262 -5072
rect -210 -5038 -144 -5022
rect -210 -5072 -194 -5038
rect -160 -5072 -144 -5038
rect -210 -5088 -144 -5072
rect -92 -5038 -26 -5022
rect -92 -5072 -76 -5038
rect -42 -5072 -26 -5038
rect -92 -5088 -26 -5072
rect 26 -5038 92 -5022
rect 26 -5072 42 -5038
rect 76 -5072 92 -5038
rect 26 -5088 92 -5072
rect 144 -5038 210 -5022
rect 144 -5072 160 -5038
rect 194 -5072 210 -5038
rect 144 -5088 210 -5072
rect 262 -5038 328 -5022
rect 262 -5072 278 -5038
rect 312 -5072 328 -5038
rect 262 -5088 328 -5072
rect 380 -5038 446 -5022
rect 380 -5072 396 -5038
rect 430 -5072 446 -5038
rect 380 -5088 446 -5072
rect 498 -5038 564 -5022
rect 498 -5072 514 -5038
rect 548 -5072 564 -5038
rect 498 -5088 564 -5072
<< polycont >>
rect -548 5038 -514 5072
rect -430 5038 -396 5072
rect -312 5038 -278 5072
rect -194 5038 -160 5072
rect -76 5038 -42 5072
rect 42 5038 76 5072
rect 160 5038 194 5072
rect 278 5038 312 5072
rect 396 5038 430 5072
rect 514 5038 548 5072
rect -548 -5072 -514 -5038
rect -430 -5072 -396 -5038
rect -312 -5072 -278 -5038
rect -194 -5072 -160 -5038
rect -76 -5072 -42 -5038
rect 42 -5072 76 -5038
rect 160 -5072 194 -5038
rect 278 -5072 312 -5038
rect 396 -5072 430 -5038
rect 514 -5072 548 -5038
<< locali >>
rect -721 5140 -625 5174
rect 625 5140 721 5174
rect -721 5078 -687 5140
rect 687 5078 721 5140
rect -564 5038 -548 5072
rect -514 5038 -498 5072
rect -446 5038 -430 5072
rect -396 5038 -380 5072
rect -328 5038 -312 5072
rect -278 5038 -262 5072
rect -210 5038 -194 5072
rect -160 5038 -144 5072
rect -92 5038 -76 5072
rect -42 5038 -26 5072
rect 26 5038 42 5072
rect 76 5038 92 5072
rect 144 5038 160 5072
rect 194 5038 210 5072
rect 262 5038 278 5072
rect 312 5038 328 5072
rect 380 5038 396 5072
rect 430 5038 446 5072
rect 498 5038 514 5072
rect 548 5038 564 5072
rect -607 4988 -573 5004
rect -607 -5004 -573 -4988
rect -489 4988 -455 5004
rect -489 -5004 -455 -4988
rect -371 4988 -337 5004
rect -371 -5004 -337 -4988
rect -253 4988 -219 5004
rect -253 -5004 -219 -4988
rect -135 4988 -101 5004
rect -135 -5004 -101 -4988
rect -17 4988 17 5004
rect -17 -5004 17 -4988
rect 101 4988 135 5004
rect 101 -5004 135 -4988
rect 219 4988 253 5004
rect 219 -5004 253 -4988
rect 337 4988 371 5004
rect 337 -5004 371 -4988
rect 455 4988 489 5004
rect 455 -5004 489 -4988
rect 573 4988 607 5004
rect 573 -5004 607 -4988
rect -564 -5072 -548 -5038
rect -514 -5072 -498 -5038
rect -446 -5072 -430 -5038
rect -396 -5072 -380 -5038
rect -328 -5072 -312 -5038
rect -278 -5072 -262 -5038
rect -210 -5072 -194 -5038
rect -160 -5072 -144 -5038
rect -92 -5072 -76 -5038
rect -42 -5072 -26 -5038
rect 26 -5072 42 -5038
rect 76 -5072 92 -5038
rect 144 -5072 160 -5038
rect 194 -5072 210 -5038
rect 262 -5072 278 -5038
rect 312 -5072 328 -5038
rect 380 -5072 396 -5038
rect 430 -5072 446 -5038
rect 498 -5072 514 -5038
rect 548 -5072 564 -5038
rect -721 -5140 -687 -5078
rect 687 -5140 721 -5078
rect -721 -5174 -625 -5140
rect 625 -5174 721 -5140
<< viali >>
rect -548 5038 -514 5072
rect -430 5038 -396 5072
rect -312 5038 -278 5072
rect -194 5038 -160 5072
rect -76 5038 -42 5072
rect 42 5038 76 5072
rect 160 5038 194 5072
rect 278 5038 312 5072
rect 396 5038 430 5072
rect 514 5038 548 5072
rect -607 -4988 -573 4988
rect -489 -4988 -455 4988
rect -371 -4988 -337 4988
rect -253 -4988 -219 4988
rect -135 -4988 -101 4988
rect -17 -4988 17 4988
rect 101 -4988 135 4988
rect 219 -4988 253 4988
rect 337 -4988 371 4988
rect 455 -4988 489 4988
rect 573 -4988 607 4988
rect -548 -5072 -514 -5038
rect -430 -5072 -396 -5038
rect -312 -5072 -278 -5038
rect -194 -5072 -160 -5038
rect -76 -5072 -42 -5038
rect 42 -5072 76 -5038
rect 160 -5072 194 -5038
rect 278 -5072 312 -5038
rect 396 -5072 430 -5038
rect 514 -5072 548 -5038
<< metal1 >>
rect -560 5072 -502 5078
rect -560 5038 -548 5072
rect -514 5038 -502 5072
rect -560 5032 -502 5038
rect -442 5072 -384 5078
rect -442 5038 -430 5072
rect -396 5038 -384 5072
rect -442 5032 -384 5038
rect -324 5072 -266 5078
rect -324 5038 -312 5072
rect -278 5038 -266 5072
rect -324 5032 -266 5038
rect -206 5072 -148 5078
rect -206 5038 -194 5072
rect -160 5038 -148 5072
rect -206 5032 -148 5038
rect -88 5072 -30 5078
rect -88 5038 -76 5072
rect -42 5038 -30 5072
rect -88 5032 -30 5038
rect 30 5072 88 5078
rect 30 5038 42 5072
rect 76 5038 88 5072
rect 30 5032 88 5038
rect 148 5072 206 5078
rect 148 5038 160 5072
rect 194 5038 206 5072
rect 148 5032 206 5038
rect 266 5072 324 5078
rect 266 5038 278 5072
rect 312 5038 324 5072
rect 266 5032 324 5038
rect 384 5072 442 5078
rect 384 5038 396 5072
rect 430 5038 442 5072
rect 384 5032 442 5038
rect 502 5072 560 5078
rect 502 5038 514 5072
rect 548 5038 560 5072
rect 502 5032 560 5038
rect -613 4988 -567 5000
rect -613 -4988 -607 4988
rect -573 -4988 -567 4988
rect -613 -5000 -567 -4988
rect -495 4988 -449 5000
rect -495 -4988 -489 4988
rect -455 -4988 -449 4988
rect -495 -5000 -449 -4988
rect -377 4988 -331 5000
rect -377 -4988 -371 4988
rect -337 -4988 -331 4988
rect -377 -5000 -331 -4988
rect -259 4988 -213 5000
rect -259 -4988 -253 4988
rect -219 -4988 -213 4988
rect -259 -5000 -213 -4988
rect -141 4988 -95 5000
rect -141 -4988 -135 4988
rect -101 -4988 -95 4988
rect -141 -5000 -95 -4988
rect -23 4988 23 5000
rect -23 -4988 -17 4988
rect 17 -4988 23 4988
rect -23 -5000 23 -4988
rect 95 4988 141 5000
rect 95 -4988 101 4988
rect 135 -4988 141 4988
rect 95 -5000 141 -4988
rect 213 4988 259 5000
rect 213 -4988 219 4988
rect 253 -4988 259 4988
rect 213 -5000 259 -4988
rect 331 4988 377 5000
rect 331 -4988 337 4988
rect 371 -4988 377 4988
rect 331 -5000 377 -4988
rect 449 4988 495 5000
rect 449 -4988 455 4988
rect 489 -4988 495 4988
rect 449 -5000 495 -4988
rect 567 4988 613 5000
rect 567 -4988 573 4988
rect 607 -4988 613 4988
rect 567 -5000 613 -4988
rect -560 -5038 -502 -5032
rect -560 -5072 -548 -5038
rect -514 -5072 -502 -5038
rect -560 -5078 -502 -5072
rect -442 -5038 -384 -5032
rect -442 -5072 -430 -5038
rect -396 -5072 -384 -5038
rect -442 -5078 -384 -5072
rect -324 -5038 -266 -5032
rect -324 -5072 -312 -5038
rect -278 -5072 -266 -5038
rect -324 -5078 -266 -5072
rect -206 -5038 -148 -5032
rect -206 -5072 -194 -5038
rect -160 -5072 -148 -5038
rect -206 -5078 -148 -5072
rect -88 -5038 -30 -5032
rect -88 -5072 -76 -5038
rect -42 -5072 -30 -5038
rect -88 -5078 -30 -5072
rect 30 -5038 88 -5032
rect 30 -5072 42 -5038
rect 76 -5072 88 -5038
rect 30 -5078 88 -5072
rect 148 -5038 206 -5032
rect 148 -5072 160 -5038
rect 194 -5072 206 -5038
rect 148 -5078 206 -5072
rect 266 -5038 324 -5032
rect 266 -5072 278 -5038
rect 312 -5072 324 -5038
rect 266 -5078 324 -5072
rect 384 -5038 442 -5032
rect 384 -5072 396 -5038
rect 430 -5072 442 -5038
rect 384 -5078 442 -5072
rect 502 -5038 560 -5032
rect 502 -5072 514 -5038
rect 548 -5072 560 -5038
rect 502 -5078 560 -5072
<< properties >>
string FIXED_BBOX -704 -5157 704 5157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 50 l 0.300 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
