** sch_path: /home/harsh/design/xschem/cs_amplifier.sch
.subckt cs_amplifier vdd output input gnd
*.PININFO input:I vdd:B gnd:B output:O
XM1 output input gnd gnd sky130_fd_pr__nfet_01v8 L=0.30 W=50 nf=10 m=1
XR1 output vdd gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.175 mult=1 m=1
.ends
.end
