* NGSPICE file created from pfd.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N a_1462_47#
+ a_543_47# a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289#
+ a_1108_47# a_1217_47# a_1659_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 Q_N a_1659_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.155 ps=1.31 w=1 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR a_1283_21# a_1659_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1522 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 VGND a_1283_21# a_1659_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 VPWR a_1659_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X18 VGND a_1659_47# Q_N VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X20 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X21 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X26 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10025 ps=0.985 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X29 Q_N a_1659_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1522 ps=1.335 w=1 l=0.15
X31 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X32 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X33 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X34 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
C0 a_1217_47# a_761_289# 4.2e-19
C1 RESET_B a_1462_47# 0.002879f
C2 Q_N a_193_47# 9.35e-20
C3 a_193_47# a_27_47# 0.906454f
C4 VPWR D 0.081188f
C5 a_193_47# a_1270_413# 1.46e-19
C6 Q RESET_B 8.5e-19
C7 a_1283_21# a_761_289# 3.17e-21
C8 Q_N VPB 0.004225f
C9 a_27_47# VPB 0.261873f
C10 VPWR a_651_413# 0.12856f
C11 Q a_193_47# 1.19e-19
C12 a_1108_47# VPWR 0.171084f
C13 VGND a_761_289# 0.073384f
C14 Q VPB 0.002023f
C15 Q_N a_27_47# 1.53e-20
C16 a_1283_21# D 2.77e-22
C17 VPWR CLK 0.017406f
C18 a_1108_47# a_1217_47# 0.007416f
C19 Q_N Q 0.0061f
C20 Q a_27_47# 3.03e-20
C21 a_1108_47# a_1283_21# 0.245854f
C22 a_639_47# a_761_289# 3.16e-19
C23 VGND D 0.051614f
C24 RESET_B a_761_289# 0.166114f
C25 a_543_47# a_761_289# 0.209641f
C26 VPWR a_1283_21# 0.156931f
C27 a_193_47# a_761_289# 0.186387f
C28 a_1108_47# VGND 0.147486f
C29 a_448_47# D 0.155634f
C30 a_1108_47# a_1659_47# 0.00277f
C31 RESET_B D 4.72e-19
C32 a_543_47# D 7.35e-20
C33 VPB a_761_289# 0.099418f
C34 VPWR VGND 0.096782f
C35 CLK VGND 0.017208f
C36 a_193_47# D 0.217945f
C37 a_1659_47# VPWR 0.205837f
C38 a_651_413# RESET_B 0.012196f
C39 a_543_47# a_651_413# 0.057222f
C40 a_1108_47# RESET_B 0.236601f
C41 a_543_47# a_1108_47# 7.99e-20
C42 a_27_47# a_761_289# 0.07009f
C43 a_805_47# a_761_289# 3.69e-19
C44 a_1270_413# a_761_289# 2.6e-19
C45 a_1217_47# VGND 9.68e-19
C46 a_193_47# a_651_413# 0.034619f
C47 D VPB 0.137565f
C48 a_448_47# VPWR 0.068142f
C49 a_1108_47# a_193_47# 0.125324f
C50 VPWR RESET_B 0.065186f
C51 a_543_47# VPWR 0.100285f
C52 CLK RESET_B 1.09e-19
C53 a_1283_21# VGND 0.2208f
C54 a_651_413# VPB 0.013543f
C55 a_1659_47# a_1283_21# 0.303605f
C56 a_27_47# D 0.132849f
C57 a_1108_47# VPB 0.111392f
C58 a_193_47# VPWR 0.395736f
C59 a_193_47# CLK 7.94e-19
C60 a_1217_47# RESET_B 6.03e-19
C61 a_651_413# a_27_47# 9.73e-19
C62 VPWR VPB 0.250676f
C63 a_448_47# a_1283_21# 1.11e-21
C64 CLK VPB 0.069345f
C65 Q_N a_1108_47# 1.34e-19
C66 a_1108_47# a_27_47# 0.102355f
C67 a_1283_21# RESET_B 0.277236f
C68 a_543_47# a_1283_21# 3.83e-21
C69 a_1217_47# a_193_47# 2.36e-20
C70 a_1108_47# a_1270_413# 0.006453f
C71 a_1659_47# VGND 0.13852f
C72 a_193_47# a_1283_21# 0.042424f
C73 Q_N VPWR 0.157089f
C74 VPWR a_27_47# 0.152295f
C75 a_27_47# CLK 0.233602f
C76 a_639_47# VGND 0.008634f
C77 VPWR a_1270_413# 7.19e-19
C78 a_448_47# VGND 0.0661f
C79 VGND RESET_B 0.28755f
C80 a_543_47# VGND 0.122935f
C81 a_1283_21# VPB 0.2414f
C82 Q VPWR 0.014118f
C83 a_1659_47# RESET_B 0.00263f
C84 a_1217_47# a_27_47# 2.56e-19
C85 a_193_47# VGND 0.063057f
C86 a_639_47# a_448_47# 4.61e-19
C87 a_639_47# RESET_B 9.54e-19
C88 a_1659_47# a_193_47# 6.89e-19
C89 Q_N a_1283_21# 0.002658f
C90 a_1283_21# a_27_47# 0.043643f
C91 a_543_47# a_639_47# 0.013793f
C92 a_448_47# RESET_B 2.45e-19
C93 a_543_47# a_448_47# 0.049827f
C94 VGND VPB 0.013806f
C95 a_543_47# RESET_B 0.153272f
C96 a_1283_21# a_1462_47# 0.007399f
C97 a_639_47# a_193_47# 2.28e-19
C98 a_1659_47# VPB 0.073099f
C99 a_448_47# a_193_47# 0.064178f
C100 Q a_1283_21# 0.053245f
C101 a_193_47# RESET_B 0.026903f
C102 a_543_47# a_193_47# 0.229804f
C103 a_651_413# a_761_289# 0.097745f
C104 Q_N VGND 0.142765f
C105 a_27_47# VGND 0.253971f
C106 a_805_47# VGND 0.00579f
C107 a_1108_47# a_761_289# 0.051162f
C108 a_448_47# VPB 0.014137f
C109 Q_N a_1659_47# 0.145144f
C110 a_1659_47# a_27_47# 5.63e-20
C111 RESET_B VPB 0.138482f
C112 VGND a_1462_47# 0.002121f
C113 a_543_47# VPB 0.095793f
C114 Q VGND 0.114874f
C115 VPWR a_761_289# 0.10497f
C116 a_639_47# a_27_47# 0.001881f
C117 a_193_47# VPB 0.170861f
C118 a_448_47# a_27_47# 0.093133f
C119 Q a_1659_47# 0.185134f
C120 Q_N RESET_B 2.83e-19
C121 a_27_47# RESET_B 0.296336f
C122 a_805_47# RESET_B 0.003155f
C123 a_543_47# a_27_47# 0.115353f
C124 a_543_47# a_805_47# 0.001705f
C125 a_1270_413# RESET_B 2.06e-19
C126 Q_N VNB 0.025191f
C127 Q VNB 0.003804f
C128 VGND VNB 1.24553f
C129 VPWR VNB 1.02447f
C130 RESET_B VNB 0.260034f
C131 D VNB 0.159894f
C132 CLK VNB 0.195254f
C133 VPB VNB 2.19949f
C134 a_1659_47# VNB 0.21348f
C135 a_651_413# VNB 0.004694f
C136 a_448_47# VNB 0.013901f
C137 a_1108_47# VNB 0.127984f
C138 a_1283_21# VNB 0.492394f
C139 a_543_47# VNB 0.157869f
C140 a_761_289# VNB 0.120848f
C141 a_193_47# VNB 0.272482f
C142 a_27_47# VNB 0.495595f
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X a_147_75# a_61_75#
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
C0 a_61_75# a_147_75# 0.006569f
C1 B X 0.002798f
C2 VGND VPB 0.009503f
C3 VGND a_61_75# 0.125003f
C4 A X 1.84e-19
C5 VPB a_61_75# 0.087048f
C6 B A 0.096585f
C7 VPWR a_147_75# 6.31e-19
C8 VGND VPWR 0.07134f
C9 VPB VPWR 0.090199f
C10 a_61_75# VPWR 0.158516f
C11 a_147_75# X 5.82e-19
C12 VGND X 0.153129f
C13 VPB X 0.005513f
C14 a_61_75# X 0.149596f
C15 B VGND 0.011526f
C16 B VPB 0.064248f
C17 B a_61_75# 0.142002f
C18 A VGND 0.015556f
C19 A VPB 0.08239f
C20 A a_61_75# 0.085863f
C21 VPWR X 0.194597f
C22 B VPWR 0.012524f
C23 A VPWR 0.040281f
C24 VGND a_147_75# 0.004769f
C25 VGND VNB 0.390327f
C26 X VNB 0.027496f
C27 B VNB 0.111386f
C28 A VNB 0.177011f
C29 VPWR VNB 0.349659f
C30 VPB VNB 0.604764f
C31 a_61_75# VNB 0.263837f
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
C0 A VPWR 0.098226f
C1 VGND VPB 0.006668f
C2 Y VPWR 0.361779f
C3 A Y 0.359887f
C4 VPWR VPB 0.065385f
C5 A VPB 0.141975f
C6 VGND VPWR 0.050092f
C7 A VGND 0.081909f
C8 Y VPB 0.015896f
C9 VGND Y 0.262586f
C10 VGND VNB 0.326816f
C11 Y VNB 0.084947f
C12 VPWR VNB 0.296394f
C13 A VNB 0.451855f
C14 VPB VNB 0.516168f
.ends

.subckt pfd VSS VDD A QA QB B
Xx1 A VDD x4/Y VSS VSS VDD VDD QA x1/Q_N x1/a_1462_47# x1/a_543_47# x1/a_651_413#
+ x1/a_193_47# x1/a_805_47# x1/a_448_47# x1/a_639_47# x1/a_1283_21# x1/a_761_289#
+ x1/a_1108_47# x1/a_1217_47# x1/a_1659_47# x1/a_1270_413# x1/a_27_47# sky130_fd_sc_hd__dfrbp_2
Xx2 QA QB VSS VSS VDD VDD x4/A x2/a_147_75# x2/a_61_75# sky130_fd_sc_hd__and2_2
Xx3 B VDD x4/Y VSS VSS VDD VDD QB x3/Q_N x3/a_1462_47# x3/a_543_47# x3/a_651_413#
+ x3/a_193_47# x3/a_805_47# x3/a_448_47# x3/a_639_47# x3/a_1283_21# x3/a_761_289#
+ x3/a_1108_47# x3/a_1217_47# x3/a_1659_47# x3/a_1270_413# x3/a_27_47# sky130_fd_sc_hd__dfrbp_2
Xx4 x4/A VSS VSS VDD VDD x4/Y sky130_fd_sc_hd__inv_4
C0 x3/a_27_47# B 0.043337f
C1 x4/Y x1/a_805_47# 0.001305f
C2 VDD x2/a_147_75# -1.11e-19
C3 A x4/Y 0.002095f
C4 QB x3/a_1283_21# 0.027088f
C5 VSS x2/a_61_75# 0.020248f
C6 x3/a_27_47# x1/a_27_47# 0.001178f
C7 x3/a_543_47# x1/a_761_289# 1.16e-21
C8 x4/A x3/a_193_47# 0.003466f
C9 VSS x3/a_805_47# 5.87e-20
C10 VDD x2/a_61_75# 0.009586f
C11 x1/a_27_47# x1/a_193_47# 1.14e-31
C12 QA VSS 0.244183f
C13 x1/a_27_47# x1/Q_N -4.19e-21
C14 x1/a_27_47# B 2.18e-20
C15 x3/a_1283_21# x3/a_27_47# -1.93e-20
C16 x3/a_27_47# x1/a_448_47# 2.34e-21
C17 A x1/a_543_47# 7.41e-19
C18 x3/a_1108_47# VSS 0.001492f
C19 VSS x3/a_1659_47# 0.006969f
C20 VDD QA 0.248217f
C21 VSS x3/a_1217_47# 4.21e-20
C22 A x1/a_761_289# 1.68e-19
C23 x3/a_1283_21# B 2.73e-20
C24 VDD x1/a_1217_47# 3.04e-20
C25 VSS x1/a_1283_21# -2.42e-19
C26 QB x3/a_193_47# 0.001069f
C27 x3/a_1108_47# VDD 6.45e-19
C28 VDD x3/a_1659_47# 0.001758f
C29 VSS x4/A 0.07421f
C30 QB x3/a_448_47# 1.46e-21
C31 x4/Y x2/a_61_75# 0.001599f
C32 VDD x1/a_1283_21# 0.012573f
C33 VSS x3/a_1270_413# 2.14e-20
C34 x4/Y x3/a_805_47# 2.28e-19
C35 x1/a_1659_47# x2/a_61_75# 3.18e-19
C36 x3/a_1283_21# x1/a_1108_47# 5.52e-21
C37 VDD x4/A 0.097844f
C38 QA x4/Y 0.04045f
C39 VDD x3/a_1270_413# 2.27e-20
C40 QA x3/Q_N 2.73e-19
C41 x3/a_193_47# x1/a_193_47# 2.32e-20
C42 x4/Y x1/a_1217_47# 2.31e-19
C43 x3/a_193_47# B 0.001688f
C44 QA x1/a_1659_47# 0.042064f
C45 x3/a_1108_47# x4/Y 0.006025f
C46 x4/Y x3/a_1659_47# 0.001136f
C47 QB VSS 0.415471f
C48 x3/a_761_289# x4/A 3.7e-19
C49 x4/Y x3/a_1217_47# 3.38e-20
C50 VDD x1/a_639_47# 4.12e-19
C51 x3/a_448_47# B 4.84e-19
C52 x4/Y x1/a_1283_21# 0.001536f
C53 x1/a_1659_47# x3/a_1659_47# 6.03e-19
C54 VDD QB 0.21605f
C55 x1/a_1283_21# x1/a_1659_47# -5.68e-32
C56 x4/Y x4/A 0.034848f
C57 QA x1/a_543_47# 5.19e-19
C58 x3/a_27_47# VSS -3.34e-19
C59 x1/a_27_47# x3/a_193_47# 9.04e-19
C60 x4/Y x3/a_1270_413# 1.2e-19
C61 QA x1/a_761_289# 4.1e-19
C62 x3/a_761_289# QB 8.51e-19
C63 x1/a_27_47# x3/a_448_47# 1.46e-21
C64 x3/a_1462_47# B 1.32e-20
C65 VSS B 0.01686f
C66 VDD x3/a_27_47# 0.002338f
C67 x4/Y x1/a_639_47# 0.001727f
C68 x3/a_193_47# x1/a_448_47# 2.22e-21
C69 VDD x1/a_193_47# 0.028809f
C70 VDD x1/Q_N 8.46e-19
C71 VDD B 0.029871f
C72 QB x4/Y 0.050099f
C73 x4/A x1/a_543_47# 0.003818f
C74 QB x3/Q_N 0.031307f
C75 x4/A x1/a_761_289# 4.33e-19
C76 QB x1/a_1659_47# 0.00212f
C77 x1/a_27_47# VSS -9.91e-19
C78 x3/a_651_413# QB 1.34e-19
C79 VSS x1/a_1108_47# 9.07e-20
C80 x3/a_543_47# x4/A 0.004131f
C81 x3/a_761_289# x1/a_193_47# 7.83e-22
C82 x3/a_761_289# B 2.15e-19
C83 x3/a_27_47# x4/Y 0.049203f
C84 x3/a_27_47# x3/Q_N -4.19e-21
C85 VDD x1/a_27_47# 0.049247f
C86 A x1/a_1283_21# 1.92e-19
C87 x3/a_1283_21# VSS 0.003083f
C88 VDD x1/a_1108_47# 0.001433f
C89 x4/Y x1/a_193_47# 0.003487f
C90 x4/Y x1/Q_N 1.16e-19
C91 B x3/a_639_47# 9.63e-20
C92 x4/Y B 0.005244f
C93 QA x2/a_147_75# 2e-19
C94 VDD x3/a_1283_21# 8.33e-19
C95 VDD x1/a_448_47# 0.003631f
C96 x3/a_761_289# x1/a_27_47# 2.37e-21
C97 QB x3/a_543_47# 4.01e-19
C98 VDD x1/a_651_413# 0.001301f
C99 x3/a_27_47# x1/a_543_47# 7.98e-21
C100 x3/a_27_47# x1/a_761_289# 2.74e-22
C101 x1/a_27_47# x4/Y 0.00875f
C102 x4/Y x1/a_1108_47# 0.003351f
C103 QA x2/a_61_75# 0.017342f
C104 VSS x3/a_193_47# 0.002595f
C105 x3/a_761_289# x1/a_651_413# 1.45e-21
C106 x1/a_27_47# x1/a_1659_47# -2.46e-20
C107 VDD x1/a_1462_47# 4.58e-20
C108 x2/a_61_75# x3/a_1659_47# 3.86e-19
C109 x3/a_543_47# x1/a_193_47# 2.29e-20
C110 x3/a_1283_21# x4/Y 0.003988f
C111 x4/Y x1/a_448_47# 0.001434f
C112 x3/a_543_47# B 3.89e-19
C113 VDD x3/a_193_47# 0.019344f
C114 x1/a_1283_21# x2/a_61_75# 0.004166f
C115 QA x1/a_1217_47# 1.11e-19
C116 x3/a_1283_21# x1/a_1659_47# 2.55e-20
C117 x1/a_651_413# x4/Y 6.75e-19
C118 x3/a_27_47# A 2.71e-19
C119 QA x3/a_1659_47# 0.001696f
C120 VDD x3/a_448_47# 0.002796f
C121 x4/A x2/a_61_75# 0.008941f
C122 QA x1/a_1283_21# 0.024967f
C123 QB x2/a_147_75# 0.001671f
C124 A x1/a_193_47# 0.001839f
C125 A B 0.005041f
C126 x1/a_27_47# x3/a_543_47# 1.4e-20
C127 VSS x3/a_1462_47# 1.39e-19
C128 x1/a_1462_47# x4/Y 2.93e-19
C129 x3/a_1108_47# x1/a_1283_21# 4.12e-20
C130 QA x4/A 0.007719f
C131 x1/a_1283_21# x3/a_1659_47# 3.88e-20
C132 x4/Y x3/a_193_47# 0.052946f
C133 VDD VSS 1.387443f
C134 x3/a_1108_47# x4/A 3.44e-19
C135 QB x2/a_61_75# 0.044533f
C136 x3/a_448_47# x4/Y 0.00253f
C137 A x1/a_27_47# 0.042843f
C138 A x1/a_1108_47# 1.35e-19
C139 x4/A x1/a_1283_21# 5.22e-19
C140 x3/a_761_289# VSS 8.85e-19
C141 QB QA 0.04773f
C142 A x1/a_448_47# 5.3e-19
C143 x3/a_193_47# x1/a_543_47# 2.55e-21
C144 x3/a_1108_47# QB 0.003904f
C145 x3/a_761_289# VDD 0.001132f
C146 QB x3/a_1659_47# 0.056973f
C147 x4/Y x3/a_1462_47# 1.45e-20
C148 VSS x3/a_639_47# 2.72e-20
C149 x3/a_193_47# x1/a_761_289# 3.27e-21
C150 VSS x4/Y 0.21309f
C151 VSS x3/Q_N 0.003831f
C152 QB x1/a_1283_21# 2.57e-19
C153 VSS x1/a_1659_47# 7.05e-19
C154 x3/a_651_413# VSS 5.67e-20
C155 VDD x4/Y 0.369261f
C156 B x3/a_805_47# 3.53e-20
C157 QB x4/A 0.015612f
C158 VDD x3/Q_N 2.66e-32
C159 x3/a_27_47# x3/a_1659_47# -2.46e-20
C160 QA x1/a_193_47# 4.04e-19
C161 QA x1/Q_N 0.027754f
C162 QB x3/a_1270_413# 6.91e-20
C163 VDD x1/a_1659_47# 0.006558f
C164 x3/a_651_413# VDD 0.001256f
C165 x1/Q_N x3/a_1659_47# 2.35e-20
C166 x3/a_1108_47# B 6.22e-20
C167 x3/a_761_289# x4/Y 0.017561f
C168 VSS x1/a_543_47# 1.11e-34
C169 B x3/a_1217_47# 1.9e-20
C170 x3/a_27_47# x4/A 0.002202f
C171 VSS x1/a_761_289# 1.18e-19
C172 x3/a_543_47# VSS 8.55e-19
C173 QA x1/a_27_47# 0.001354f
C174 x3/a_1283_21# x2/a_61_75# 0.004423f
C175 VDD x1/a_543_47# 0.006327f
C176 QA x1/a_1108_47# 0.002246f
C177 x4/Y x3/a_639_47# 1.03e-19
C178 x4/A x1/a_193_47# 0.00332f
C179 x4/Y x3/Q_N 5.99e-20
C180 VDD x1/a_761_289# 0.003739f
C181 VDD x3/a_543_47# 0.002217f
C182 x3/a_1108_47# x1/a_1108_47# 5.91e-19
C183 x4/Y x1/a_1659_47# -2e-20
C184 x3/a_1283_21# QA 1.43e-19
C185 x3/Q_N x1/a_1659_47# 4.61e-20
C186 x3/a_651_413# x4/Y 0.010022f
C187 QA x1/a_448_47# 2.27e-20
C188 x3/a_761_289# x1/a_543_47# 4.39e-21
C189 x1/a_27_47# x1/a_1283_21# -1.12e-20
C190 A VSS 0.019504f
C191 QB x3/a_27_47# 7.99e-19
C192 x3/a_761_289# x1/a_761_289# 5.95e-19
C193 x3/a_1283_21# x3/a_1659_47# 5.68e-32
C194 VDD x1/a_805_47# 1.61e-19
C195 x1/a_27_47# x4/A 0.003279f
C196 VDD x1/a_1270_413# 2.63e-20
C197 x4/A x1/a_1108_47# 3.36e-19
C198 QB x1/Q_N 2.45e-19
C199 VDD A 0.303684f
C200 x4/Y x1/a_543_47# 0.006791f
C201 x3/a_1283_21# x1/a_1283_21# 0.002542f
C202 x4/Y x1/a_761_289# 0.006611f
C203 QA x1/a_1462_47# 3.2e-19
C204 x3/a_543_47# x4/Y 0.016593f
C205 x3/a_1283_21# x4/A 6.39e-19
C206 VSS x2/a_147_75# 5.7e-19
C207 x3/a_651_413# x1/a_761_289# 6.52e-21
C208 x3/a_27_47# x1/a_193_47# 7.46e-19
C209 VSS 0 2.91701f
C210 x4/Y 0 0.934107f
C211 x4/A 0 0.533512f
C212 VDD 0 8.719146f
C213 x3/Q_N 0 0.025191f
C214 QB 0 0.66652f
C215 B 0 0.37907f
C216 x3/a_1659_47# 0 0.21348f
C217 x3/a_651_413# 0 0.004694f
C218 x3/a_448_47# 0 0.013901f
C219 x3/a_1108_47# 0 0.127984f
C220 x3/a_1283_21# 0 0.492394f
C221 x3/a_543_47# 0 0.157869f
C222 x3/a_761_289# 0 0.120848f
C223 x3/a_193_47# 0 0.272482f
C224 x3/a_27_47# 0 0.495595f
C225 QA 0 0.658428f
C226 x2/a_61_75# 0 0.263837f
C227 x1/Q_N 0 0.025191f
C228 A 0 0.493384f
C229 x1/a_1659_47# 0 0.21348f
C230 x1/a_651_413# 0 0.004694f
C231 x1/a_448_47# 0 0.013901f
C232 x1/a_1108_47# 0 0.127984f
C233 x1/a_1283_21# 0 0.492394f
C234 x1/a_543_47# 0 0.157869f
C235 x1/a_761_289# 0 0.120848f
C236 x1/a_193_47# 0 0.272482f
C237 x1/a_27_47# 0 0.495595f
.ends

