magic
tech sky130A
magscale 1 2
timestamp 1706843384
<< error_s >>
rect 608 2380 610 2450
<< locali >>
rect 114 1876 206 2312
<< viali >>
rect 704 576 920 624
<< metal1 >>
rect 382 2380 392 2462
rect 542 2380 552 2462
rect 1334 2452 1534 2522
rect 920 2388 930 2448
rect 1040 2388 1050 2448
rect 1334 2386 1368 2452
rect 1500 2386 1534 2452
rect 1334 2322 1534 2386
rect -354 2100 -154 2156
rect -354 2006 -312 2100
rect -210 2006 -154 2100
rect -354 1956 -154 2006
rect -328 1844 -16 1846
rect 106 1844 406 1850
rect -328 1788 406 1844
rect -420 1588 -220 1788
rect -168 1786 406 1788
rect 528 1786 1280 1850
rect -328 728 -218 1588
rect 74 1562 84 1730
rect 144 1562 154 1730
rect 308 1566 318 1734
rect 378 1566 388 1734
rect 546 1568 556 1736
rect 616 1568 626 1736
rect 784 1568 794 1736
rect 854 1568 864 1736
rect 1020 1570 1030 1738
rect 1090 1570 1100 1738
rect 1258 1572 1268 1740
rect 1328 1572 1338 1740
rect 194 804 204 972
rect 264 804 274 972
rect 432 806 442 974
rect 502 806 512 974
rect 662 810 672 978
rect 732 810 742 978
rect 898 810 908 978
rect 968 810 978 978
rect 1134 800 1144 968
rect 1204 800 1214 968
rect -328 726 112 728
rect -328 674 1274 726
rect -328 664 112 674
rect 692 624 744 630
rect 886 624 932 630
rect 692 576 704 624
rect 920 576 932 624
rect 692 570 744 576
rect 734 568 744 570
rect 886 570 932 576
rect 886 568 896 570
rect 728 418 928 476
rect 728 336 778 418
rect 870 336 928 418
rect 728 276 928 336
<< via1 >>
rect 392 2380 542 2462
rect 930 2388 1040 2448
rect 1368 2386 1500 2452
rect -312 2006 -210 2100
rect 84 1562 144 1730
rect 318 1566 378 1734
rect 556 1568 616 1736
rect 794 1568 854 1736
rect 1030 1570 1090 1738
rect 1268 1572 1328 1740
rect 204 804 264 972
rect 442 806 502 974
rect 672 810 732 978
rect 908 810 968 978
rect 1144 800 1204 968
rect 744 624 886 630
rect 744 576 886 624
rect 744 568 886 576
rect 778 336 870 418
<< metal2 >>
rect 392 2462 542 2472
rect 392 2370 542 2380
rect 930 2450 1040 2458
rect 1368 2452 1500 2462
rect 930 2448 1368 2450
rect 1040 2390 1368 2448
rect 930 2378 1040 2388
rect 1500 2390 1536 2450
rect 1368 2376 1500 2386
rect 406 2124 528 2370
rect -326 2100 528 2124
rect -326 2006 -312 2100
rect -210 2006 528 2100
rect -326 1994 528 2006
rect 84 1732 144 1740
rect 318 1734 378 1744
rect 60 1730 318 1732
rect 60 1576 84 1730
rect 144 1576 318 1730
rect 84 1552 144 1562
rect 406 1732 528 1994
rect 556 1736 616 1746
rect 378 1576 556 1732
rect 318 1556 378 1566
rect 794 1736 854 1746
rect 616 1578 794 1732
rect 616 1576 688 1578
rect 746 1576 794 1578
rect 556 1558 616 1568
rect 1030 1738 1090 1748
rect 854 1576 1030 1732
rect 794 1558 854 1568
rect 1268 1740 1328 1750
rect 1090 1576 1268 1732
rect 1030 1560 1090 1570
rect 1328 1576 1352 1732
rect 1268 1562 1328 1572
rect 442 982 502 984
rect 672 982 732 988
rect 908 982 968 988
rect 184 978 1220 982
rect 184 974 672 978
rect 184 972 442 974
rect 184 804 204 972
rect 264 806 442 972
rect 502 810 672 974
rect 732 810 908 978
rect 968 968 1220 978
rect 968 810 1144 968
rect 502 806 1144 810
rect 264 804 1144 806
rect 184 800 1144 804
rect 1204 800 1220 968
rect 184 798 1220 800
rect 204 794 264 798
rect 442 796 502 798
rect 760 640 868 798
rect 1144 790 1204 798
rect 744 630 886 640
rect 744 558 886 568
rect 760 428 868 558
rect 760 418 870 428
rect 760 336 778 418
rect 760 326 870 336
rect 760 320 868 326
use sky130_fd_pr__nfet_01v8_4H4H2H  XM1
timestamp 1706794580
transform 1 0 704 0 1 1257
box -757 -710 757 710
use sky130_fd_pr__res_xhigh_po_0p35_4SYHMP  XR1
timestamp 1706691097
transform 0 1 574 -1 0 2415
box -201 -632 201 632
<< labels >>
flabel metal1 -420 1588 -220 1788 0 FreeSans 256 0 0 0 input
port 2 nsew
flabel metal1 728 276 928 476 0 FreeSans 256 0 0 0 gnd
port 3 nsew
flabel metal1 -354 1956 -154 2156 0 FreeSans 256 0 0 0 output
port 1 nsew
flabel metal1 1334 2322 1534 2522 0 FreeSans 256 0 0 0 vdd
port 0 nsew
<< end >>
