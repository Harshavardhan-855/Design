magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< error_p >>
rect -407 114 -349 120
rect -191 114 -133 120
rect 25 114 83 120
rect 241 114 299 120
rect 457 114 515 120
rect -407 80 -395 114
rect -191 80 -179 114
rect 25 80 37 114
rect 241 80 253 114
rect 457 80 469 114
rect -407 74 -349 80
rect -191 74 -133 80
rect 25 74 83 80
rect 241 74 299 80
rect 457 74 515 80
rect -515 -80 -457 -74
rect -299 -80 -241 -74
rect -83 -80 -25 -74
rect 133 -80 191 -74
rect 349 -80 407 -74
rect -515 -114 -503 -80
rect -299 -114 -287 -80
rect -83 -114 -71 -80
rect 133 -114 145 -80
rect 349 -114 361 -80
rect -515 -120 -457 -114
rect -299 -120 -241 -114
rect -83 -120 -25 -114
rect 133 -120 191 -114
rect 349 -120 407 -114
<< pwell >>
rect -707 -252 707 252
<< nmos >>
rect -511 -42 -461 42
rect -403 -42 -353 42
rect -295 -42 -245 42
rect -187 -42 -137 42
rect -79 -42 -29 42
rect 29 -42 79 42
rect 137 -42 187 42
rect 245 -42 295 42
rect 353 -42 403 42
rect 461 -42 511 42
<< ndiff >>
rect -569 30 -511 42
rect -569 -30 -557 30
rect -523 -30 -511 30
rect -569 -42 -511 -30
rect -461 30 -403 42
rect -461 -30 -449 30
rect -415 -30 -403 30
rect -461 -42 -403 -30
rect -353 30 -295 42
rect -353 -30 -341 30
rect -307 -30 -295 30
rect -353 -42 -295 -30
rect -245 30 -187 42
rect -245 -30 -233 30
rect -199 -30 -187 30
rect -245 -42 -187 -30
rect -137 30 -79 42
rect -137 -30 -125 30
rect -91 -30 -79 30
rect -137 -42 -79 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 79 30 137 42
rect 79 -30 91 30
rect 125 -30 137 30
rect 79 -42 137 -30
rect 187 30 245 42
rect 187 -30 199 30
rect 233 -30 245 30
rect 187 -42 245 -30
rect 295 30 353 42
rect 295 -30 307 30
rect 341 -30 353 30
rect 295 -42 353 -30
rect 403 30 461 42
rect 403 -30 415 30
rect 449 -30 461 30
rect 403 -42 461 -30
rect 511 30 569 42
rect 511 -30 523 30
rect 557 -30 569 30
rect 511 -42 569 -30
<< ndiffc >>
rect -557 -30 -523 30
rect -449 -30 -415 30
rect -341 -30 -307 30
rect -233 -30 -199 30
rect -125 -30 -91 30
rect -17 -30 17 30
rect 91 -30 125 30
rect 199 -30 233 30
rect 307 -30 341 30
rect 415 -30 449 30
rect 523 -30 557 30
<< psubdiff >>
rect -671 182 -575 216
rect 575 182 671 216
rect -671 120 -637 182
rect 637 120 671 182
rect -671 -182 -637 -120
rect 637 -182 671 -120
rect -671 -216 -575 -182
rect 575 -216 671 -182
<< psubdiffcont >>
rect -575 182 575 216
rect -671 -120 -637 120
rect 637 -120 671 120
rect -575 -216 575 -182
<< poly >>
rect -411 114 -345 130
rect -411 80 -395 114
rect -361 80 -345 114
rect -511 42 -461 68
rect -411 64 -345 80
rect -195 114 -129 130
rect -195 80 -179 114
rect -145 80 -129 114
rect -403 42 -353 64
rect -295 42 -245 68
rect -195 64 -129 80
rect 21 114 87 130
rect 21 80 37 114
rect 71 80 87 114
rect -187 42 -137 64
rect -79 42 -29 68
rect 21 64 87 80
rect 237 114 303 130
rect 237 80 253 114
rect 287 80 303 114
rect 29 42 79 64
rect 137 42 187 68
rect 237 64 303 80
rect 453 114 519 130
rect 453 80 469 114
rect 503 80 519 114
rect 245 42 295 64
rect 353 42 403 68
rect 453 64 519 80
rect 461 42 511 64
rect -511 -64 -461 -42
rect -519 -80 -453 -64
rect -403 -68 -353 -42
rect -295 -64 -245 -42
rect -519 -114 -503 -80
rect -469 -114 -453 -80
rect -519 -130 -453 -114
rect -303 -80 -237 -64
rect -187 -68 -137 -42
rect -79 -64 -29 -42
rect -303 -114 -287 -80
rect -253 -114 -237 -80
rect -303 -130 -237 -114
rect -87 -80 -21 -64
rect 29 -68 79 -42
rect 137 -64 187 -42
rect -87 -114 -71 -80
rect -37 -114 -21 -80
rect -87 -130 -21 -114
rect 129 -80 195 -64
rect 245 -68 295 -42
rect 353 -64 403 -42
rect 129 -114 145 -80
rect 179 -114 195 -80
rect 129 -130 195 -114
rect 345 -80 411 -64
rect 461 -68 511 -42
rect 345 -114 361 -80
rect 395 -114 411 -80
rect 345 -130 411 -114
<< polycont >>
rect -395 80 -361 114
rect -179 80 -145 114
rect 37 80 71 114
rect 253 80 287 114
rect 469 80 503 114
rect -503 -114 -469 -80
rect -287 -114 -253 -80
rect -71 -114 -37 -80
rect 145 -114 179 -80
rect 361 -114 395 -80
<< locali >>
rect -671 182 -575 216
rect 575 182 671 216
rect -671 120 -637 182
rect 637 120 671 182
rect -411 80 -395 114
rect -361 80 -345 114
rect -195 80 -179 114
rect -145 80 -129 114
rect 21 80 37 114
rect 71 80 87 114
rect 237 80 253 114
rect 287 80 303 114
rect 453 80 469 114
rect 503 80 519 114
rect -557 30 -523 46
rect -557 -46 -523 -30
rect -449 30 -415 46
rect -449 -46 -415 -30
rect -341 30 -307 46
rect -341 -46 -307 -30
rect -233 30 -199 46
rect -233 -46 -199 -30
rect -125 30 -91 46
rect -125 -46 -91 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 91 30 125 46
rect 91 -46 125 -30
rect 199 30 233 46
rect 199 -46 233 -30
rect 307 30 341 46
rect 307 -46 341 -30
rect 415 30 449 46
rect 415 -46 449 -30
rect 523 30 557 46
rect 523 -46 557 -30
rect -519 -114 -503 -80
rect -469 -114 -453 -80
rect -303 -114 -287 -80
rect -253 -114 -237 -80
rect -87 -114 -71 -80
rect -37 -114 -21 -80
rect 129 -114 145 -80
rect 179 -114 195 -80
rect 345 -114 361 -80
rect 395 -114 411 -80
rect -671 -182 -637 -120
rect 637 -182 671 -120
rect -671 -216 -575 -182
rect 575 -216 671 -182
<< viali >>
rect -395 80 -361 114
rect -179 80 -145 114
rect 37 80 71 114
rect 253 80 287 114
rect 469 80 503 114
rect -557 -30 -523 30
rect -449 -30 -415 30
rect -341 -30 -307 30
rect -233 -30 -199 30
rect -125 -30 -91 30
rect -17 -30 17 30
rect 91 -30 125 30
rect 199 -30 233 30
rect 307 -30 341 30
rect 415 -30 449 30
rect 523 -30 557 30
rect -503 -114 -469 -80
rect -287 -114 -253 -80
rect -71 -114 -37 -80
rect 145 -114 179 -80
rect 361 -114 395 -80
<< metal1 >>
rect -407 114 -349 120
rect -407 80 -395 114
rect -361 80 -349 114
rect -407 74 -349 80
rect -191 114 -133 120
rect -191 80 -179 114
rect -145 80 -133 114
rect -191 74 -133 80
rect 25 114 83 120
rect 25 80 37 114
rect 71 80 83 114
rect 25 74 83 80
rect 241 114 299 120
rect 241 80 253 114
rect 287 80 299 114
rect 241 74 299 80
rect 457 114 515 120
rect 457 80 469 114
rect 503 80 515 114
rect 457 74 515 80
rect -563 30 -517 42
rect -563 -30 -557 30
rect -523 -30 -517 30
rect -563 -42 -517 -30
rect -455 30 -409 42
rect -455 -30 -449 30
rect -415 -30 -409 30
rect -455 -42 -409 -30
rect -347 30 -301 42
rect -347 -30 -341 30
rect -307 -30 -301 30
rect -347 -42 -301 -30
rect -239 30 -193 42
rect -239 -30 -233 30
rect -199 -30 -193 30
rect -239 -42 -193 -30
rect -131 30 -85 42
rect -131 -30 -125 30
rect -91 -30 -85 30
rect -131 -42 -85 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 85 30 131 42
rect 85 -30 91 30
rect 125 -30 131 30
rect 85 -42 131 -30
rect 193 30 239 42
rect 193 -30 199 30
rect 233 -30 239 30
rect 193 -42 239 -30
rect 301 30 347 42
rect 301 -30 307 30
rect 341 -30 347 30
rect 301 -42 347 -30
rect 409 30 455 42
rect 409 -30 415 30
rect 449 -30 455 30
rect 409 -42 455 -30
rect 517 30 563 42
rect 517 -30 523 30
rect 557 -30 563 30
rect 517 -42 563 -30
rect -515 -80 -457 -74
rect -515 -114 -503 -80
rect -469 -114 -457 -80
rect -515 -120 -457 -114
rect -299 -80 -241 -74
rect -299 -114 -287 -80
rect -253 -114 -241 -80
rect -299 -120 -241 -114
rect -83 -80 -25 -74
rect -83 -114 -71 -80
rect -37 -114 -25 -80
rect -83 -120 -25 -114
rect 133 -80 191 -74
rect 133 -114 145 -80
rect 179 -114 191 -80
rect 133 -120 191 -114
rect 349 -80 407 -74
rect 349 -114 361 -80
rect 395 -114 407 -80
rect 349 -120 407 -114
<< properties >>
string FIXED_BBOX -654 -199 654 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.250 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
