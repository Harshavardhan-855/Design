magic
tech sky130A
magscale 1 2
timestamp 1706788245
<< pwell >>
rect -5158 -471 5158 471
<< ndiff >>
rect -5000 301 5000 313
rect -5000 267 -4988 301
rect 4988 267 5000 301
rect -5000 210 5000 267
rect -5000 -267 5000 -210
rect -5000 -301 -4988 -267
rect 4988 -301 5000 -267
rect -5000 -313 5000 -301
<< ndiffc >>
rect -4988 267 4988 301
rect -4988 -301 4988 -267
<< psubdiff >>
rect -5122 401 -5026 435
rect 5026 401 5122 435
rect -5122 339 -5088 401
rect 5088 339 5122 401
rect -5122 -401 -5088 -339
rect 5088 -401 5122 -339
rect -5122 -435 -5026 -401
rect 5026 -435 5122 -401
<< psubdiffcont >>
rect -5026 401 5026 435
rect -5122 -339 -5088 339
rect 5088 -339 5122 339
rect -5026 -435 5026 -401
<< ndiffres >>
rect -5000 -210 5000 210
<< locali >>
rect -5122 401 -5026 435
rect 5026 401 5122 435
rect -5122 339 -5088 401
rect 5088 339 5122 401
rect -5004 267 -4988 301
rect 4988 267 5004 301
rect -5004 -301 -4988 -267
rect 4988 -301 5004 -267
rect -5122 -401 -5088 -339
rect 5088 -401 5122 -339
rect -5122 -435 -5026 -401
rect 5026 -435 5122 -401
<< viali >>
rect -4988 267 4988 301
rect -4988 227 4988 267
rect -4988 -267 4988 -227
rect -4988 -301 4988 -267
<< metal1 >>
rect -5000 301 5000 307
rect -5000 227 -4988 301
rect 4988 227 5000 301
rect -5000 221 5000 227
rect -5000 -227 5000 -221
rect -5000 -301 -4988 -227
rect 4988 -301 5000 -227
rect -5000 -307 5000 -301
<< properties >>
string FIXED_BBOX -5105 -418 5105 418
string gencell sky130_fd_pr__res_generic_nd
string library sky130
string parameters w 50 l 2.10 m 1 nx 1 wmin 0.42 lmin 2.10 rho 120 val 5.045 dummy 0 dw 0.05 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
