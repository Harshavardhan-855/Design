magic
tech sky130A
magscale 1 2
timestamp 1709903010
<< error_s >>
rect 3374 -562 4324 -516
rect 3374 -568 3396 -562
rect 4214 -816 4324 -562
rect 3314 -1353 3372 -1347
rect 3314 -1387 3326 -1353
rect 3314 -1393 3372 -1387
rect 3522 -1396 3524 -1330
rect 3550 -1353 3608 -1347
rect 3550 -1387 3562 -1353
rect 3550 -1393 3608 -1387
rect 3351 -1626 3370 -1426
rect 3379 -1654 3398 -1434
rect 5680 -1454 5700 -1422
rect 3528 -1586 3543 -1470
rect 3735 -1486 3769 -1468
rect 5708 -1482 5728 -1450
rect 3556 -1558 3571 -1498
rect 3735 -1522 3805 -1486
rect 5101 -1512 5159 -1506
rect 5219 -1512 5277 -1506
rect 5337 -1512 5395 -1506
rect 5455 -1512 5513 -1506
rect 5573 -1512 5631 -1506
rect 3752 -1556 3823 -1522
rect 4251 -1556 4286 -1522
rect 4822 -1539 4856 -1521
rect 3314 -1881 3372 -1875
rect 3432 -1881 3490 -1875
rect 3550 -1881 3608 -1875
rect 3314 -1915 3326 -1881
rect 3432 -1915 3444 -1881
rect 3550 -1915 3562 -1881
rect 3314 -1921 3372 -1915
rect 3432 -1921 3490 -1915
rect 3550 -1921 3608 -1915
rect 3752 -2017 3822 -1556
rect 4252 -1575 4286 -1556
rect 3949 -1624 4007 -1618
rect 4067 -1624 4125 -1618
rect 3949 -1658 3961 -1624
rect 4067 -1658 4079 -1624
rect 3949 -1664 4007 -1658
rect 4067 -1664 4125 -1658
rect 3949 -1934 4007 -1928
rect 4067 -1934 4125 -1928
rect 3949 -1968 3961 -1934
rect 4067 -1968 4079 -1934
rect 3949 -1974 4007 -1968
rect 4067 -1974 4125 -1968
rect 3752 -2053 3805 -2017
rect 4271 -2070 4286 -1575
rect 4305 -1609 4340 -1575
rect 4305 -2070 4339 -1609
rect 4466 -1677 4524 -1671
rect 4466 -1711 4478 -1677
rect 4466 -1717 4524 -1711
rect 4466 -1987 4524 -1981
rect 4584 -1987 4642 -1981
rect 4466 -2021 4478 -1987
rect 4584 -2021 4596 -1987
rect 4466 -2027 4524 -2021
rect 4584 -2027 4642 -2021
rect 4305 -2104 4320 -2070
rect 4786 -2123 4856 -1539
rect 5101 -1546 5113 -1512
rect 5219 -1546 5231 -1512
rect 5337 -1546 5349 -1512
rect 5455 -1546 5467 -1512
rect 5573 -1546 5585 -1512
rect 5950 -1523 6200 -1202
rect 6646 -1522 6696 -1426
rect 5101 -1552 5159 -1546
rect 5219 -1552 5277 -1546
rect 5337 -1552 5395 -1546
rect 5455 -1552 5513 -1546
rect 5573 -1552 5631 -1546
rect 5138 -1680 5148 -1642
rect 5172 -1714 5182 -1608
rect 5526 -1852 5560 -1605
rect 5680 -1678 5684 -1593
rect 5708 -1650 5712 -1572
rect 6646 -1680 6648 -1654
rect 6292 -1687 6646 -1680
rect 5876 -1705 5910 -1687
rect 5876 -1741 5946 -1705
rect 6025 -1737 6077 -1687
rect 6107 -1707 6161 -1687
rect 6101 -1733 6167 -1707
rect 6107 -1737 6161 -1733
rect 6191 -1737 6245 -1687
rect 6275 -1707 6646 -1687
rect 6269 -1716 6646 -1707
rect 6648 -1716 6674 -1680
rect 6269 -1733 6648 -1716
rect 6275 -1737 6648 -1733
rect 6292 -1741 6648 -1737
rect 5893 -1775 5964 -1741
rect 6025 -1750 6648 -1741
rect 7013 -1750 7048 -1733
rect 6025 -1762 6646 -1750
rect 6067 -1767 6201 -1762
rect 6235 -1763 6646 -1762
rect 6235 -1767 6362 -1763
rect 6369 -1767 6396 -1763
rect 6432 -1766 6646 -1763
rect 5526 -1904 5600 -1852
rect 5526 -1981 5560 -1904
rect 4983 -2040 5041 -2034
rect 5101 -2040 5159 -2034
rect 5219 -2040 5277 -2034
rect 5337 -2040 5395 -2034
rect 5455 -2040 5513 -2034
rect 5573 -2040 5631 -2034
rect 5691 -2040 5749 -2034
rect 4983 -2074 4995 -2040
rect 5101 -2074 5113 -2040
rect 5219 -2074 5231 -2040
rect 5337 -2074 5349 -2040
rect 5455 -2074 5467 -2040
rect 5573 -2074 5585 -2040
rect 5691 -2074 5703 -2040
rect 4983 -2080 5041 -2074
rect 5101 -2080 5159 -2074
rect 5219 -2080 5277 -2074
rect 5337 -2080 5395 -2074
rect 5455 -2080 5513 -2074
rect 5573 -2080 5631 -2074
rect 5691 -2080 5749 -2074
rect 4786 -2159 4839 -2123
rect 5893 -2176 5963 -1775
rect 5988 -1801 5997 -1775
rect 6292 -1784 6369 -1767
rect 6419 -1771 6646 -1766
rect 6648 -1771 6674 -1750
rect 6419 -1784 6674 -1771
rect 6062 -1832 6120 -1809
rect 6090 -1860 6120 -1837
rect 6090 -2093 6148 -2087
rect 6090 -2127 6102 -2093
rect 6090 -2133 6148 -2127
rect 5893 -2212 5946 -2176
rect 6292 -2229 6362 -1784
rect 6432 -1802 6674 -1784
rect 7014 -1751 7048 -1750
rect 7014 -1787 7084 -1751
rect 6432 -1824 6648 -1802
rect 6486 -1826 6648 -1824
rect 7031 -1821 7102 -1787
rect 6292 -2265 6345 -2229
rect 7031 -2282 7101 -1821
rect 7031 -2318 7084 -2282
rect 8370 -2371 8423 -1751
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use pfd  x1
timestamp 1708936645
transform 1 0 -786 0 1 -120
box 786 -1880 3956 334
use cp_schem  x2
timestamp 1709901343
transform 1 0 850 0 1 -984
box 2267 -1440 8916 1562
use inverter  x3
timestamp 1709276979
transform 1 0 5988 0 1 -2384
box -280 384 1040 1362
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 cp_bias
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 cp_out
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 B
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
