magic
tech sky130A
magscale 1 2
timestamp 1708425308
<< error_p >>
rect -29 1599 29 1605
rect -29 1565 -17 1599
rect -29 1559 29 1565
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -1565 29 -1559
rect -29 -1599 -17 -1565
rect -29 -1605 29 -1599
<< nwell >>
rect -226 -1737 226 1737
<< pmos >>
rect -30 118 30 1518
rect -30 -1518 30 -118
<< pdiff >>
rect -88 1506 -30 1518
rect -88 130 -76 1506
rect -42 130 -30 1506
rect -88 118 -30 130
rect 30 1506 88 1518
rect 30 130 42 1506
rect 76 130 88 1506
rect 30 118 88 130
rect -88 -130 -30 -118
rect -88 -1506 -76 -130
rect -42 -1506 -30 -130
rect -88 -1518 -30 -1506
rect 30 -130 88 -118
rect 30 -1506 42 -130
rect 76 -1506 88 -130
rect 30 -1518 88 -1506
<< pdiffc >>
rect -76 130 -42 1506
rect 42 130 76 1506
rect -76 -1506 -42 -130
rect 42 -1506 76 -130
<< nsubdiff >>
rect -190 1667 -94 1701
rect 94 1667 190 1701
rect -190 1605 -156 1667
rect 156 1605 190 1667
rect -190 -1667 -156 -1605
rect 156 -1667 190 -1605
rect -190 -1701 -94 -1667
rect 94 -1701 190 -1667
<< nsubdiffcont >>
rect -94 1667 94 1701
rect -190 -1605 -156 1605
rect 156 -1605 190 1605
rect -94 -1701 94 -1667
<< poly >>
rect -33 1599 33 1615
rect -33 1565 -17 1599
rect 17 1565 33 1599
rect -33 1549 33 1565
rect -30 1518 30 1549
rect -30 87 30 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -118 30 -87
rect -30 -1549 30 -1518
rect -33 -1565 33 -1549
rect -33 -1599 -17 -1565
rect 17 -1599 33 -1565
rect -33 -1615 33 -1599
<< polycont >>
rect -17 1565 17 1599
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -1599 17 -1565
<< locali >>
rect -190 1667 -94 1701
rect 94 1667 190 1701
rect -190 1605 -156 1667
rect 156 1605 190 1667
rect -33 1565 -17 1599
rect 17 1565 33 1599
rect -76 1506 -42 1522
rect -76 114 -42 130
rect 42 1506 76 1522
rect 42 114 76 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -130 -42 -114
rect -76 -1522 -42 -1506
rect 42 -130 76 -114
rect 42 -1522 76 -1506
rect -33 -1599 -17 -1565
rect 17 -1599 33 -1565
rect -190 -1667 -156 -1605
rect 156 -1667 190 -1605
rect -190 -1701 -94 -1667
rect 94 -1701 190 -1667
<< viali >>
rect -17 1565 17 1599
rect -76 130 -42 1506
rect 42 130 76 1506
rect -17 37 17 71
rect -17 -71 17 -37
rect -76 -1506 -42 -130
rect 42 -1506 76 -130
rect -17 -1599 17 -1565
<< metal1 >>
rect -29 1599 29 1605
rect -29 1565 -17 1599
rect 17 1565 29 1599
rect -29 1559 29 1565
rect -82 1506 -36 1518
rect -82 130 -76 1506
rect -42 130 -36 1506
rect -82 118 -36 130
rect 36 1506 82 1518
rect 36 130 42 1506
rect 76 130 82 1506
rect 36 118 82 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -130 -36 -118
rect -82 -1506 -76 -130
rect -42 -1506 -36 -130
rect -82 -1518 -36 -1506
rect 36 -130 82 -118
rect 36 -1506 42 -130
rect 76 -1506 82 -130
rect 36 -1518 82 -1506
rect -29 -1565 29 -1559
rect -29 -1599 -17 -1565
rect 17 -1599 29 -1565
rect -29 -1605 29 -1599
<< properties >>
string FIXED_BBOX -173 -1684 173 1684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 0.3 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
