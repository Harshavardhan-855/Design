magic
tech sky130A
magscale 1 2
timestamp 1709276637
<< nwell >>
rect 3344 284 3378 286
rect 3344 244 3364 284
rect 3394 8 3614 334
rect 3394 -16 3612 8
rect 1830 -458 2002 -438
rect 1830 -734 1990 -458
rect 3344 -528 3536 -486
rect 1841 -735 1990 -734
rect 1952 -744 1990 -735
rect 3416 -792 3536 -528
rect 3416 -793 3529 -792
rect 3384 -1250 3552 -1230
rect 3398 -1266 3552 -1250
rect 3342 -1302 3552 -1266
rect 3398 -1526 3552 -1302
rect 3398 -1527 3533 -1526
rect 3398 -1528 3420 -1527
<< pwell >>
rect 3346 -270 3544 -86
rect 3344 -306 3544 -270
rect 3346 -336 3544 -306
rect 2026 -874 2060 -838
rect 1876 -1092 2086 -874
rect 3370 -906 3528 -858
rect 3370 -1104 3530 -906
rect 3352 -1810 3508 -1680
rect 3300 -1880 3510 -1810
<< psubdiff >>
rect 3420 -168 3512 -144
rect 3420 -334 3512 -310
rect 1888 -906 1980 -882
rect 1888 -1072 1980 -1048
rect 3426 -936 3518 -912
rect 3426 -1102 3518 -1078
rect 3404 -1706 3496 -1682
rect 3404 -1872 3496 -1848
<< nsubdiff >>
rect 3474 246 3551 280
rect 3517 220 3551 246
rect 3517 92 3551 118
rect 3474 58 3551 92
rect 1875 -511 1952 -477
rect 1875 -537 1909 -511
rect 3418 -569 3495 -535
rect 1875 -665 1909 -639
rect 3461 -595 3495 -569
rect 1875 -699 1952 -665
rect 3461 -723 3495 -697
rect 3418 -757 3495 -723
rect 3422 -1303 3499 -1269
rect 3465 -1329 3499 -1303
rect 3465 -1457 3499 -1431
rect 3422 -1491 3499 -1457
<< psubdiffcont >>
rect 3420 -310 3512 -168
rect 1888 -1048 1980 -906
rect 3426 -1078 3518 -936
rect 3404 -1848 3496 -1706
<< nsubdiffcont >>
rect 3517 118 3551 220
rect 1875 -639 1909 -537
rect 3461 -697 3495 -595
rect 3465 -1431 3499 -1329
<< locali >>
rect 3344 284 3378 286
rect 3344 280 3504 284
rect 3344 246 3551 280
rect 3344 244 3364 246
rect 3517 220 3551 246
rect 3517 92 3551 118
rect 3474 58 3551 92
rect 1230 -82 1238 -30
rect 3420 -168 3512 -152
rect 3344 -306 3420 -272
rect 3420 -326 3512 -310
rect 1896 -462 1958 -460
rect 1896 -477 2036 -462
rect 1875 -510 2036 -477
rect 1875 -511 1938 -510
rect 1875 -537 1909 -511
rect 3358 -535 3452 -506
rect 3358 -542 3495 -535
rect 3418 -569 3495 -542
rect 1875 -665 1909 -639
rect 3461 -595 3495 -569
rect 1875 -699 1952 -665
rect 3461 -723 3495 -697
rect 1926 -776 2076 -750
rect 3418 -757 3495 -723
rect 1926 -824 1970 -776
rect 2024 -824 2076 -776
rect 2650 -780 2698 -778
rect 2392 -804 2698 -780
rect 2392 -808 2740 -804
rect 2392 -818 2984 -808
rect 1926 -846 2076 -824
rect 2654 -846 2984 -818
rect 1888 -906 1980 -890
rect 3426 -936 3518 -920
rect 1980 -1048 2030 -1024
rect 1888 -1060 2030 -1048
rect 1888 -1064 1980 -1060
rect 3360 -1078 3426 -1050
rect 3360 -1084 3518 -1078
rect 3426 -1094 3518 -1084
rect 3346 -1269 3452 -1266
rect 3346 -1302 3499 -1269
rect 3422 -1303 3499 -1302
rect 3465 -1329 3499 -1303
rect 3465 -1457 3499 -1431
rect 3422 -1491 3499 -1457
rect 3404 -1706 3496 -1690
rect 3322 -1848 3404 -1822
rect 3322 -1864 3496 -1848
<< viali >>
rect 1456 148 1492 192
rect 1180 -82 1230 -30
rect 3012 -76 3064 -34
rect 3312 -762 3348 -728
rect 1970 -824 2024 -776
rect 3122 -852 3170 -800
rect 1444 -1400 1484 -1358
rect 1168 -1624 1230 -1566
rect 3004 -1620 3052 -1572
<< metal1 >>
rect 982 242 1234 306
rect 982 106 1182 242
rect 1448 192 1498 250
rect 1448 148 1456 192
rect 1492 148 1498 192
rect 1448 130 1498 148
rect 786 -24 986 42
rect 786 -86 862 -24
rect 950 -86 986 -24
rect 786 -158 986 -86
rect 1016 -462 1104 106
rect 3638 -22 3838 20
rect 1132 -90 1142 -24
rect 1242 -90 1252 -24
rect 3002 -28 3012 -24
rect 3000 -82 3012 -28
rect 3064 -28 3074 -24
rect 3002 -86 3012 -82
rect 3064 -82 3076 -28
rect 3064 -86 3074 -82
rect 3638 -92 3700 -22
rect 3774 -92 3838 -22
rect 2007 -153 2017 -93
rect 2071 -153 2081 -93
rect 3638 -180 3838 -92
rect 3292 -336 3714 -240
rect 1018 -548 2082 -462
rect 2390 -544 2910 -450
rect 1640 -1314 1712 -548
rect 1946 -828 1956 -766
rect 2034 -828 2044 -766
rect 3290 -772 3300 -716
rect 3364 -772 3374 -716
rect 3116 -800 3176 -788
rect 3116 -806 3122 -800
rect 3170 -806 3176 -800
rect 1958 -830 2036 -828
rect 3100 -862 3110 -806
rect 3182 -862 3192 -806
rect 3116 -864 3176 -862
rect 2422 -1108 2906 -994
rect 3624 -1022 3714 -336
rect 3290 -1112 3714 -1022
rect 1431 -1358 1496 -1314
rect 1431 -1400 1444 -1358
rect 1484 -1400 1496 -1358
rect 1431 -1413 1496 -1400
rect 872 -1572 1072 -1518
rect 1156 -1566 1242 -1560
rect 1156 -1572 1168 -1566
rect 872 -1624 1168 -1572
rect 1230 -1624 1242 -1566
rect 872 -1718 1072 -1624
rect 1156 -1630 1242 -1624
rect 2972 -1628 2982 -1564
rect 3072 -1628 3082 -1564
rect 1992 -1694 2002 -1634
rect 2056 -1694 2066 -1634
rect 3624 -1674 3714 -1112
rect 3514 -1784 3714 -1674
rect 3756 -1526 3956 -1476
rect 3756 -1630 3804 -1526
rect 3890 -1630 3956 -1526
rect 3756 -1676 3956 -1630
rect 3282 -1874 3714 -1784
<< via1 >>
rect 862 -86 950 -24
rect 1142 -30 1242 -24
rect 1142 -82 1180 -30
rect 1180 -82 1230 -30
rect 1230 -82 1242 -30
rect 1142 -90 1242 -82
rect 3012 -34 3064 -24
rect 3012 -76 3064 -34
rect 3012 -86 3064 -76
rect 3700 -92 3774 -22
rect 2017 -153 2071 -93
rect 1956 -776 2034 -766
rect 1956 -824 1970 -776
rect 1970 -824 2024 -776
rect 2024 -824 2034 -776
rect 1956 -828 2034 -824
rect 3300 -728 3364 -716
rect 3300 -762 3312 -728
rect 3312 -762 3348 -728
rect 3348 -762 3364 -728
rect 3300 -772 3364 -762
rect 3110 -852 3122 -806
rect 3122 -852 3170 -806
rect 3170 -852 3182 -806
rect 3110 -862 3182 -852
rect 2982 -1572 3072 -1564
rect 2982 -1620 3004 -1572
rect 3004 -1620 3052 -1572
rect 3052 -1620 3072 -1572
rect 2982 -1628 3072 -1620
rect 2002 -1694 2056 -1634
rect 3804 -1630 3890 -1526
<< metal2 >>
rect 860 -10 1242 -8
rect 860 -22 1244 -10
rect 3012 -22 3064 -14
rect 3292 -16 3370 -14
rect 3700 -16 3774 -12
rect 3292 -22 3774 -16
rect 860 -24 1246 -22
rect 860 -86 862 -24
rect 950 -86 1142 -24
rect 860 -90 1142 -86
rect 1242 -90 1246 -24
rect 3010 -24 3700 -22
rect 3010 -76 3012 -24
rect 860 -94 1246 -90
rect 2017 -93 2071 -83
rect 860 -98 1242 -94
rect 1142 -100 1242 -98
rect 3064 -76 3700 -24
rect 3012 -96 3064 -86
rect 3292 -90 3700 -76
rect 2017 -163 2071 -153
rect 2018 -756 2068 -163
rect 1956 -766 2068 -756
rect 2034 -826 2068 -766
rect 3292 -716 3370 -90
rect 3700 -102 3774 -92
rect 3292 -770 3300 -716
rect 3364 -770 3370 -716
rect 3300 -782 3364 -772
rect 3110 -806 3182 -796
rect 2034 -828 2066 -826
rect 1956 -838 2066 -828
rect 2002 -1628 2066 -838
rect 3110 -872 3182 -862
rect 2982 -1562 3072 -1554
rect 3116 -1558 3182 -872
rect 3804 -1526 3890 -1516
rect 3104 -1562 3804 -1558
rect 2982 -1564 3804 -1562
rect 3072 -1614 3804 -1564
rect 3072 -1620 3182 -1614
rect 3116 -1624 3182 -1620
rect 1998 -1634 2090 -1628
rect 1998 -1694 2002 -1634
rect 2056 -1694 2090 -1634
rect 2982 -1638 3072 -1628
rect 3804 -1640 3890 -1630
rect 1998 -1698 2090 -1694
rect 2002 -1704 2056 -1698
use sky130_fd_sc_hd__dfrbp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform 1 0 1170 0 1 -288
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 3378 0 1 -1068
box -38 -48 590 592
use sky130_fd_sc_hd__dfrbp_2  x3
timestamp 1705271942
transform 1 0 1160 0 1 -1830
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 2474 0 1 -1040
box -38 -48 498 592
<< labels >>
flabel metal1 3514 -1874 3714 -1674 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 982 106 1182 306 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 786 -158 986 42 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 872 -1718 1072 -1518 0 FreeSans 256 0 0 0 B
port 5 nsew
flabel metal1 3756 -1676 3956 -1476 0 FreeSans 256 0 0 0 QB
port 4 nsew
flabel metal1 3638 -180 3838 20 0 FreeSans 256 0 0 0 QA
port 3 nsew
<< end >>
