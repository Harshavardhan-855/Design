magic
tech sky130A
magscale 1 2
timestamp 1706862968
<< pwell >>
rect -830 1614 310 1662
rect 1254 1600 2394 1648
rect 1256 490 2396 538
<< viali >>
rect 212 182 364 444
rect 1158 180 1310 442
rect 782 -1136 904 -1094
<< metal1 >>
rect 634 2592 834 2792
rect -832 2094 -822 2304
rect -624 2094 -614 2304
rect 640 2300 830 2592
rect -36 2114 1516 2300
rect 2016 2162 2026 2272
rect 2334 2162 2344 2272
rect -1602 1922 -1402 1982
rect -1602 1836 -1550 1922
rect -1456 1836 -1402 1922
rect -1602 1782 -1402 1836
rect 2728 1914 2928 1972
rect 2728 1824 2784 1914
rect 2878 1824 2928 1914
rect 2728 1772 2928 1824
rect -1174 1656 282 1662
rect -1178 1616 282 1656
rect -1592 1024 -1392 1104
rect -1178 1024 -1118 1616
rect -858 1614 282 1616
rect 1226 1644 2366 1648
rect 2616 1644 2652 1646
rect 1226 1600 2654 1644
rect 2332 1598 2654 1600
rect -920 1350 -910 1546
rect -854 1350 -844 1546
rect -678 1344 -668 1540
rect -612 1344 -602 1540
rect -446 1352 -436 1548
rect -380 1352 -370 1548
rect -208 1354 -198 1550
rect -142 1354 -132 1550
rect 28 1358 38 1554
rect 94 1358 104 1554
rect 260 1362 270 1558
rect 326 1362 336 1558
rect 1164 1330 1174 1522
rect 1254 1330 1264 1522
rect 1404 1332 1414 1524
rect 1494 1332 1504 1524
rect 1630 1336 1640 1528
rect 1720 1336 1730 1528
rect 1876 1332 1886 1524
rect 1966 1332 1976 1524
rect 2102 1328 2112 1520
rect 2192 1328 2202 1520
rect 2344 1340 2354 1532
rect 2434 1340 2444 1532
rect -1592 974 -1118 1024
rect -1592 904 -1392 974
rect -1178 548 -1118 974
rect 2616 1116 2652 1598
rect 2836 1116 3036 1204
rect 2616 1066 3036 1116
rect -800 604 -790 772
rect -734 604 -724 772
rect -560 614 -550 772
rect -488 614 -478 772
rect -328 620 -318 774
rect -258 620 -248 774
rect -94 614 -84 768
rect -24 614 -14 768
rect 146 620 156 774
rect 216 620 226 774
rect 1284 592 1294 794
rect 1362 592 1372 794
rect 1522 590 1532 792
rect 1600 590 1610 792
rect 1758 598 1768 800
rect 1836 598 1846 800
rect 2004 598 2014 800
rect 2082 598 2092 800
rect 2230 580 2240 782
rect 2308 580 2318 782
rect -864 548 276 550
rect -1178 504 276 548
rect -1154 502 276 504
rect 1228 536 2368 538
rect 2616 536 2652 1066
rect 2836 1004 3036 1066
rect -1154 500 -786 502
rect 1228 490 2662 536
rect 206 444 370 456
rect 206 182 212 444
rect 364 182 370 444
rect 206 170 370 182
rect 1152 442 1316 454
rect 1152 180 1158 442
rect 1310 180 1316 442
rect 1152 168 1316 180
rect -114 76 1380 118
rect -416 -434 -216 -366
rect -86 -434 -6 76
rect 240 70 1380 76
rect 178 -202 188 -10
rect 262 -202 272 -10
rect 416 -204 426 -12
rect 500 -204 510 -12
rect 656 -204 666 -12
rect 740 -204 750 -12
rect 890 -202 900 -10
rect 974 -202 984 -10
rect 1122 -200 1132 -8
rect 1206 -200 1216 -8
rect 1368 -198 1378 -6
rect 1452 -198 1462 -6
rect -416 -500 -6 -434
rect -416 -566 -216 -500
rect -86 -996 -6 -500
rect 292 -932 302 -740
rect 376 -932 386 -740
rect 542 -926 552 -734
rect 626 -926 636 -734
rect 774 -922 784 -730
rect 858 -922 868 -730
rect 1002 -940 1012 -748
rect 1086 -940 1096 -748
rect 1240 -942 1250 -750
rect 1324 -942 1334 -750
rect 240 -996 1380 -994
rect -86 -1036 1380 -996
rect -52 -1042 1380 -1036
rect 790 -1088 800 -1084
rect 770 -1094 800 -1088
rect 880 -1088 890 -1084
rect 880 -1094 916 -1088
rect 770 -1136 782 -1094
rect 904 -1136 916 -1094
rect 770 -1142 800 -1136
rect 790 -1152 800 -1142
rect 880 -1142 916 -1136
rect 880 -1152 890 -1142
rect 744 -1332 944 -1276
rect 744 -1420 802 -1332
rect 886 -1420 944 -1332
rect 744 -1476 944 -1420
<< via1 >>
rect -822 2094 -624 2304
rect 2026 2162 2334 2272
rect -1550 1836 -1456 1922
rect 2784 1824 2878 1914
rect -910 1350 -854 1546
rect -668 1344 -612 1540
rect -436 1352 -380 1548
rect -198 1354 -142 1550
rect 38 1358 94 1554
rect 270 1362 326 1558
rect 1174 1330 1254 1522
rect 1414 1332 1494 1524
rect 1640 1336 1720 1528
rect 1886 1332 1966 1524
rect 2112 1328 2192 1520
rect 2354 1340 2434 1532
rect -790 604 -734 772
rect -550 614 -488 772
rect -318 620 -258 774
rect -84 614 -24 768
rect 156 620 216 774
rect 1294 592 1362 794
rect 1532 590 1600 792
rect 1768 598 1836 800
rect 2014 598 2082 800
rect 2240 580 2308 782
rect 188 -202 262 -10
rect 426 -204 500 -12
rect 666 -204 740 -12
rect 900 -202 974 -10
rect 1132 -200 1206 -8
rect 1378 -198 1452 -6
rect 302 -932 376 -740
rect 552 -926 626 -734
rect 784 -922 858 -730
rect 1012 -940 1086 -748
rect 1250 -942 1324 -750
rect 800 -1094 880 -1084
rect 800 -1136 880 -1094
rect 800 -1152 880 -1136
rect 802 -1420 886 -1332
<< metal2 >>
rect -822 2304 -624 2314
rect -826 2094 -822 2302
rect 2026 2272 2334 2282
rect 2026 2152 2334 2162
rect -826 2084 -624 2094
rect -1550 1922 -1456 1932
rect -826 1914 -692 2084
rect -1456 1836 -692 1914
rect -1550 1826 -1456 1836
rect -910 1552 -854 1556
rect -826 1552 -692 1836
rect 2202 1902 2298 2152
rect 2784 1914 2878 1924
rect 2202 1826 2784 1902
rect -436 1552 -380 1558
rect -198 1552 -142 1560
rect 38 1554 94 1564
rect -926 1550 38 1552
rect -926 1548 -198 1550
rect -926 1546 -436 1548
rect -926 1364 -910 1546
rect -854 1540 -436 1546
rect -854 1364 -668 1540
rect -910 1340 -854 1350
rect -612 1364 -436 1540
rect -668 1334 -612 1344
rect -380 1364 -198 1548
rect -436 1342 -380 1352
rect -142 1364 38 1550
rect -198 1344 -142 1354
rect 270 1558 326 1568
rect 94 1364 270 1552
rect 38 1348 94 1358
rect 326 1364 338 1552
rect 2202 1540 2298 1826
rect 2784 1814 2878 1824
rect 2354 1540 2434 1542
rect 1156 1532 2452 1540
rect 1156 1528 2354 1532
rect 1156 1524 1640 1528
rect 1156 1522 1414 1524
rect 270 1352 326 1362
rect 1156 1336 1174 1522
rect 1254 1336 1414 1522
rect 1174 1320 1254 1330
rect 1494 1336 1640 1524
rect 1720 1524 2354 1528
rect 1720 1336 1886 1524
rect 1414 1322 1494 1332
rect 1640 1326 1720 1336
rect 1966 1520 2354 1524
rect 1966 1336 2112 1520
rect 1886 1322 1966 1332
rect 2192 1340 2354 1520
rect 2434 1340 2452 1532
rect 2192 1336 2452 1340
rect 2354 1330 2434 1336
rect 2112 1318 2192 1328
rect 1294 794 1362 804
rect 1532 794 1600 802
rect 1768 800 1836 810
rect -790 772 -734 782
rect -550 772 -488 782
rect -318 774 -258 784
rect -824 620 -790 772
rect -734 620 -550 772
rect -488 620 -318 772
rect -84 772 -24 778
rect 156 774 216 784
rect -258 768 156 772
rect -258 620 -84 768
rect -550 604 -488 614
rect -318 610 -258 620
rect -24 620 156 768
rect 216 730 236 772
rect 1258 730 1294 794
rect 216 632 1294 730
rect 216 620 236 632
rect -84 604 -24 614
rect 156 610 216 620
rect -790 594 -734 604
rect 188 -4 262 0
rect 426 -4 500 -2
rect 666 -4 740 -2
rect 774 -4 856 632
rect 1258 598 1294 632
rect 1362 792 1768 794
rect 1362 598 1532 792
rect 1294 582 1362 592
rect 1600 598 1768 792
rect 2014 800 2082 810
rect 1836 598 2014 794
rect 2082 782 2344 794
rect 2082 598 2240 782
rect 1532 580 1600 590
rect 1768 588 1836 598
rect 2014 588 2082 598
rect 2308 598 2344 782
rect 2240 570 2308 580
rect 900 -4 974 0
rect 1132 -4 1206 2
rect 1378 -4 1452 4
rect 164 -6 1478 -4
rect 164 -8 1378 -6
rect 164 -10 1132 -8
rect 164 -194 188 -10
rect 262 -12 900 -10
rect 262 -194 426 -12
rect 188 -212 262 -202
rect 500 -194 666 -12
rect 426 -214 500 -204
rect 740 -194 900 -12
rect 666 -214 740 -204
rect 974 -194 1132 -10
rect 900 -212 974 -202
rect 1206 -194 1378 -8
rect 1132 -210 1206 -200
rect 1452 -194 1478 -6
rect 1378 -208 1452 -198
rect 302 -732 376 -730
rect 552 -732 626 -724
rect 784 -730 858 -720
rect 274 -734 784 -732
rect 274 -740 552 -734
rect 274 -932 302 -740
rect 376 -926 552 -740
rect 626 -922 784 -734
rect 858 -748 1346 -732
rect 858 -922 1012 -748
rect 626 -926 1012 -922
rect 376 -932 1012 -926
rect 302 -942 376 -932
rect 552 -936 626 -932
rect 788 -1084 896 -932
rect 1086 -750 1346 -748
rect 1086 -932 1250 -750
rect 1012 -950 1086 -940
rect 1324 -932 1346 -750
rect 1250 -952 1324 -942
rect 788 -1152 800 -1084
rect 880 -1152 896 -1084
rect 788 -1332 896 -1152
rect 788 -1420 802 -1332
rect 886 -1420 896 -1332
rect 788 -1424 896 -1420
rect 802 -1430 886 -1424
use sky130_fd_pr__res_generic_po_XJGAA7  R1
timestamp 1706794580
transform 0 1 -240 -1 0 2206
box -266 -846 266 846
use sky130_fd_pr__res_generic_po_XJGAA7  R2
timestamp 1706794580
transform 0 -1 1710 -1 0 2220
box -266 -846 266 846
use sky130_fd_pr__nfet_01v8_4H4H2H  XM1
timestamp 1706794580
transform 1 0 -289 0 1 1082
box -757 -710 757 710
use sky130_fd_pr__nfet_01v8_4H4H2H  XM2
timestamp 1706794580
transform 1 0 1801 0 1 1066
box -757 -710 757 710
use sky130_fd_pr__nfet_01v8_4H4H2H  XM3
timestamp 1706794580
transform 1 0 817 0 1 -458
box -757 -710 757 710
<< labels >>
flabel metal1 -1592 904 -1392 1104 0 FreeSans 256 0 0 0 inp1
port 2 nsew
flabel metal1 634 2592 834 2792 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 -1602 1782 -1402 1982 0 FreeSans 256 0 0 0 out1
port 5 nsew
flabel metal1 744 -1476 944 -1276 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 2728 1772 2928 1972 0 FreeSans 256 0 0 0 out2
port 4 nsew
flabel metal1 2836 1004 3036 1204 0 FreeSans 256 0 0 0 inp2
port 3 nsew
flabel metal1 -416 -566 -216 -366 0 FreeSans 256 0 0 0 vbias
port 6 nsew
<< end >>
