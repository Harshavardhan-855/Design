magic
tech sky130A
magscale 1 2
timestamp 1707817411
<< error_p >>
rect -29 781 29 787
rect -29 747 -17 781
rect -29 741 29 747
rect -29 -747 29 -741
rect -29 -781 -17 -747
rect -29 -787 29 -781
<< nwell >>
rect -226 -919 226 919
<< pmos >>
rect -30 -700 30 700
<< pdiff >>
rect -88 688 -30 700
rect -88 -688 -76 688
rect -42 -688 -30 688
rect -88 -700 -30 -688
rect 30 688 88 700
rect 30 -688 42 688
rect 76 -688 88 688
rect 30 -700 88 -688
<< pdiffc >>
rect -76 -688 -42 688
rect 42 -688 76 688
<< nsubdiff >>
rect -190 849 -94 883
rect 94 849 190 883
rect -190 787 -156 849
rect 156 787 190 849
rect -190 -849 -156 -787
rect 156 -849 190 -787
rect -190 -883 -94 -849
rect 94 -883 190 -849
<< nsubdiffcont >>
rect -94 849 94 883
rect -190 -787 -156 787
rect 156 -787 190 787
rect -94 -883 94 -849
<< poly >>
rect -33 781 33 797
rect -33 747 -17 781
rect 17 747 33 781
rect -33 731 33 747
rect -30 700 30 731
rect -30 -731 30 -700
rect -33 -747 33 -731
rect -33 -781 -17 -747
rect 17 -781 33 -747
rect -33 -797 33 -781
<< polycont >>
rect -17 747 17 781
rect -17 -781 17 -747
<< locali >>
rect -190 849 -94 883
rect 94 849 190 883
rect -190 787 -156 849
rect 156 787 190 849
rect -33 747 -17 781
rect 17 747 33 781
rect -76 688 -42 704
rect -76 -704 -42 -688
rect 42 688 76 704
rect 42 -704 76 -688
rect -33 -781 -17 -747
rect 17 -781 33 -747
rect -190 -849 -156 -787
rect 156 -849 190 -787
rect -190 -883 -94 -849
rect 94 -883 190 -849
<< viali >>
rect -17 747 17 781
rect -76 -688 -42 688
rect 42 -688 76 688
rect -17 -781 17 -747
<< metal1 >>
rect -29 781 29 787
rect -29 747 -17 781
rect 17 747 29 781
rect -29 741 29 747
rect -82 688 -36 700
rect -82 -688 -76 688
rect -42 -688 -36 688
rect -82 -700 -36 -688
rect 36 688 82 700
rect 36 -688 42 688
rect 76 -688 82 688
rect 36 -700 82 -688
rect -29 -747 29 -741
rect -29 -781 -17 -747
rect 17 -781 29 -747
rect -29 -787 29 -781
<< properties >>
string FIXED_BBOX -173 -866 173 866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
