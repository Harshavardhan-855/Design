magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -4205 372 -4147 378
rect -4013 372 -3955 378
rect -3821 372 -3763 378
rect -3629 372 -3571 378
rect -3437 372 -3379 378
rect -3245 372 -3187 378
rect -3053 372 -2995 378
rect -2861 372 -2803 378
rect -2669 372 -2611 378
rect -2477 372 -2419 378
rect -2285 372 -2227 378
rect -2093 372 -2035 378
rect -1901 372 -1843 378
rect -1709 372 -1651 378
rect -1517 372 -1459 378
rect -1325 372 -1267 378
rect -1133 372 -1075 378
rect -941 372 -883 378
rect -749 372 -691 378
rect -557 372 -499 378
rect -365 372 -307 378
rect -173 372 -115 378
rect 19 372 77 378
rect 211 372 269 378
rect 403 372 461 378
rect 595 372 653 378
rect 787 372 845 378
rect 979 372 1037 378
rect 1171 372 1229 378
rect 1363 372 1421 378
rect 1555 372 1613 378
rect 1747 372 1805 378
rect 1939 372 1997 378
rect 2131 372 2189 378
rect 2323 372 2381 378
rect 2515 372 2573 378
rect 2707 372 2765 378
rect 2899 372 2957 378
rect 3091 372 3149 378
rect 3283 372 3341 378
rect 3475 372 3533 378
rect 3667 372 3725 378
rect 3859 372 3917 378
rect 4051 372 4109 378
rect 4243 372 4301 378
rect -4205 338 -4193 372
rect -4013 338 -4001 372
rect -3821 338 -3809 372
rect -3629 338 -3617 372
rect -3437 338 -3425 372
rect -3245 338 -3233 372
rect -3053 338 -3041 372
rect -2861 338 -2849 372
rect -2669 338 -2657 372
rect -2477 338 -2465 372
rect -2285 338 -2273 372
rect -2093 338 -2081 372
rect -1901 338 -1889 372
rect -1709 338 -1697 372
rect -1517 338 -1505 372
rect -1325 338 -1313 372
rect -1133 338 -1121 372
rect -941 338 -929 372
rect -749 338 -737 372
rect -557 338 -545 372
rect -365 338 -353 372
rect -173 338 -161 372
rect 19 338 31 372
rect 211 338 223 372
rect 403 338 415 372
rect 595 338 607 372
rect 787 338 799 372
rect 979 338 991 372
rect 1171 338 1183 372
rect 1363 338 1375 372
rect 1555 338 1567 372
rect 1747 338 1759 372
rect 1939 338 1951 372
rect 2131 338 2143 372
rect 2323 338 2335 372
rect 2515 338 2527 372
rect 2707 338 2719 372
rect 2899 338 2911 372
rect 3091 338 3103 372
rect 3283 338 3295 372
rect 3475 338 3487 372
rect 3667 338 3679 372
rect 3859 338 3871 372
rect 4051 338 4063 372
rect 4243 338 4255 372
rect -4205 332 -4147 338
rect -4013 332 -3955 338
rect -3821 332 -3763 338
rect -3629 332 -3571 338
rect -3437 332 -3379 338
rect -3245 332 -3187 338
rect -3053 332 -2995 338
rect -2861 332 -2803 338
rect -2669 332 -2611 338
rect -2477 332 -2419 338
rect -2285 332 -2227 338
rect -2093 332 -2035 338
rect -1901 332 -1843 338
rect -1709 332 -1651 338
rect -1517 332 -1459 338
rect -1325 332 -1267 338
rect -1133 332 -1075 338
rect -941 332 -883 338
rect -749 332 -691 338
rect -557 332 -499 338
rect -365 332 -307 338
rect -173 332 -115 338
rect 19 332 77 338
rect 211 332 269 338
rect 403 332 461 338
rect 595 332 653 338
rect 787 332 845 338
rect 979 332 1037 338
rect 1171 332 1229 338
rect 1363 332 1421 338
rect 1555 332 1613 338
rect 1747 332 1805 338
rect 1939 332 1997 338
rect 2131 332 2189 338
rect 2323 332 2381 338
rect 2515 332 2573 338
rect 2707 332 2765 338
rect 2899 332 2957 338
rect 3091 332 3149 338
rect 3283 332 3341 338
rect 3475 332 3533 338
rect 3667 332 3725 338
rect 3859 332 3917 338
rect 4051 332 4109 338
rect 4243 332 4301 338
rect -4301 -338 -4243 -332
rect -4109 -338 -4051 -332
rect -3917 -338 -3859 -332
rect -3725 -338 -3667 -332
rect -3533 -338 -3475 -332
rect -3341 -338 -3283 -332
rect -3149 -338 -3091 -332
rect -2957 -338 -2899 -332
rect -2765 -338 -2707 -332
rect -2573 -338 -2515 -332
rect -2381 -338 -2323 -332
rect -2189 -338 -2131 -332
rect -1997 -338 -1939 -332
rect -1805 -338 -1747 -332
rect -1613 -338 -1555 -332
rect -1421 -338 -1363 -332
rect -1229 -338 -1171 -332
rect -1037 -338 -979 -332
rect -845 -338 -787 -332
rect -653 -338 -595 -332
rect -461 -338 -403 -332
rect -269 -338 -211 -332
rect -77 -338 -19 -332
rect 115 -338 173 -332
rect 307 -338 365 -332
rect 499 -338 557 -332
rect 691 -338 749 -332
rect 883 -338 941 -332
rect 1075 -338 1133 -332
rect 1267 -338 1325 -332
rect 1459 -338 1517 -332
rect 1651 -338 1709 -332
rect 1843 -338 1901 -332
rect 2035 -338 2093 -332
rect 2227 -338 2285 -332
rect 2419 -338 2477 -332
rect 2611 -338 2669 -332
rect 2803 -338 2861 -332
rect 2995 -338 3053 -332
rect 3187 -338 3245 -332
rect 3379 -338 3437 -332
rect 3571 -338 3629 -332
rect 3763 -338 3821 -332
rect 3955 -338 4013 -332
rect 4147 -338 4205 -332
rect -4301 -372 -4289 -338
rect -4109 -372 -4097 -338
rect -3917 -372 -3905 -338
rect -3725 -372 -3713 -338
rect -3533 -372 -3521 -338
rect -3341 -372 -3329 -338
rect -3149 -372 -3137 -338
rect -2957 -372 -2945 -338
rect -2765 -372 -2753 -338
rect -2573 -372 -2561 -338
rect -2381 -372 -2369 -338
rect -2189 -372 -2177 -338
rect -1997 -372 -1985 -338
rect -1805 -372 -1793 -338
rect -1613 -372 -1601 -338
rect -1421 -372 -1409 -338
rect -1229 -372 -1217 -338
rect -1037 -372 -1025 -338
rect -845 -372 -833 -338
rect -653 -372 -641 -338
rect -461 -372 -449 -338
rect -269 -372 -257 -338
rect -77 -372 -65 -338
rect 115 -372 127 -338
rect 307 -372 319 -338
rect 499 -372 511 -338
rect 691 -372 703 -338
rect 883 -372 895 -338
rect 1075 -372 1087 -338
rect 1267 -372 1279 -338
rect 1459 -372 1471 -338
rect 1651 -372 1663 -338
rect 1843 -372 1855 -338
rect 2035 -372 2047 -338
rect 2227 -372 2239 -338
rect 2419 -372 2431 -338
rect 2611 -372 2623 -338
rect 2803 -372 2815 -338
rect 2995 -372 3007 -338
rect 3187 -372 3199 -338
rect 3379 -372 3391 -338
rect 3571 -372 3583 -338
rect 3763 -372 3775 -338
rect 3955 -372 3967 -338
rect 4147 -372 4159 -338
rect -4301 -378 -4243 -372
rect -4109 -378 -4051 -372
rect -3917 -378 -3859 -372
rect -3725 -378 -3667 -372
rect -3533 -378 -3475 -372
rect -3341 -378 -3283 -372
rect -3149 -378 -3091 -372
rect -2957 -378 -2899 -372
rect -2765 -378 -2707 -372
rect -2573 -378 -2515 -372
rect -2381 -378 -2323 -372
rect -2189 -378 -2131 -372
rect -1997 -378 -1939 -372
rect -1805 -378 -1747 -372
rect -1613 -378 -1555 -372
rect -1421 -378 -1363 -372
rect -1229 -378 -1171 -372
rect -1037 -378 -979 -372
rect -845 -378 -787 -372
rect -653 -378 -595 -372
rect -461 -378 -403 -372
rect -269 -378 -211 -372
rect -77 -378 -19 -372
rect 115 -378 173 -372
rect 307 -378 365 -372
rect 499 -378 557 -372
rect 691 -378 749 -372
rect 883 -378 941 -372
rect 1075 -378 1133 -372
rect 1267 -378 1325 -372
rect 1459 -378 1517 -372
rect 1651 -378 1709 -372
rect 1843 -378 1901 -372
rect 2035 -378 2093 -372
rect 2227 -378 2285 -372
rect 2419 -378 2477 -372
rect 2611 -378 2669 -372
rect 2803 -378 2861 -372
rect 2995 -378 3053 -372
rect 3187 -378 3245 -372
rect 3379 -378 3437 -372
rect 3571 -378 3629 -372
rect 3763 -378 3821 -372
rect 3955 -378 4013 -372
rect 4147 -378 4205 -372
<< pwell >>
rect -4487 -510 4487 510
<< nmos >>
rect -4287 -300 -4257 300
rect -4191 -300 -4161 300
rect -4095 -300 -4065 300
rect -3999 -300 -3969 300
rect -3903 -300 -3873 300
rect -3807 -300 -3777 300
rect -3711 -300 -3681 300
rect -3615 -300 -3585 300
rect -3519 -300 -3489 300
rect -3423 -300 -3393 300
rect -3327 -300 -3297 300
rect -3231 -300 -3201 300
rect -3135 -300 -3105 300
rect -3039 -300 -3009 300
rect -2943 -300 -2913 300
rect -2847 -300 -2817 300
rect -2751 -300 -2721 300
rect -2655 -300 -2625 300
rect -2559 -300 -2529 300
rect -2463 -300 -2433 300
rect -2367 -300 -2337 300
rect -2271 -300 -2241 300
rect -2175 -300 -2145 300
rect -2079 -300 -2049 300
rect -1983 -300 -1953 300
rect -1887 -300 -1857 300
rect -1791 -300 -1761 300
rect -1695 -300 -1665 300
rect -1599 -300 -1569 300
rect -1503 -300 -1473 300
rect -1407 -300 -1377 300
rect -1311 -300 -1281 300
rect -1215 -300 -1185 300
rect -1119 -300 -1089 300
rect -1023 -300 -993 300
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
rect 993 -300 1023 300
rect 1089 -300 1119 300
rect 1185 -300 1215 300
rect 1281 -300 1311 300
rect 1377 -300 1407 300
rect 1473 -300 1503 300
rect 1569 -300 1599 300
rect 1665 -300 1695 300
rect 1761 -300 1791 300
rect 1857 -300 1887 300
rect 1953 -300 1983 300
rect 2049 -300 2079 300
rect 2145 -300 2175 300
rect 2241 -300 2271 300
rect 2337 -300 2367 300
rect 2433 -300 2463 300
rect 2529 -300 2559 300
rect 2625 -300 2655 300
rect 2721 -300 2751 300
rect 2817 -300 2847 300
rect 2913 -300 2943 300
rect 3009 -300 3039 300
rect 3105 -300 3135 300
rect 3201 -300 3231 300
rect 3297 -300 3327 300
rect 3393 -300 3423 300
rect 3489 -300 3519 300
rect 3585 -300 3615 300
rect 3681 -300 3711 300
rect 3777 -300 3807 300
rect 3873 -300 3903 300
rect 3969 -300 3999 300
rect 4065 -300 4095 300
rect 4161 -300 4191 300
rect 4257 -300 4287 300
<< ndiff >>
rect -4349 288 -4287 300
rect -4349 -288 -4337 288
rect -4303 -288 -4287 288
rect -4349 -300 -4287 -288
rect -4257 288 -4191 300
rect -4257 -288 -4241 288
rect -4207 -288 -4191 288
rect -4257 -300 -4191 -288
rect -4161 288 -4095 300
rect -4161 -288 -4145 288
rect -4111 -288 -4095 288
rect -4161 -300 -4095 -288
rect -4065 288 -3999 300
rect -4065 -288 -4049 288
rect -4015 -288 -3999 288
rect -4065 -300 -3999 -288
rect -3969 288 -3903 300
rect -3969 -288 -3953 288
rect -3919 -288 -3903 288
rect -3969 -300 -3903 -288
rect -3873 288 -3807 300
rect -3873 -288 -3857 288
rect -3823 -288 -3807 288
rect -3873 -300 -3807 -288
rect -3777 288 -3711 300
rect -3777 -288 -3761 288
rect -3727 -288 -3711 288
rect -3777 -300 -3711 -288
rect -3681 288 -3615 300
rect -3681 -288 -3665 288
rect -3631 -288 -3615 288
rect -3681 -300 -3615 -288
rect -3585 288 -3519 300
rect -3585 -288 -3569 288
rect -3535 -288 -3519 288
rect -3585 -300 -3519 -288
rect -3489 288 -3423 300
rect -3489 -288 -3473 288
rect -3439 -288 -3423 288
rect -3489 -300 -3423 -288
rect -3393 288 -3327 300
rect -3393 -288 -3377 288
rect -3343 -288 -3327 288
rect -3393 -300 -3327 -288
rect -3297 288 -3231 300
rect -3297 -288 -3281 288
rect -3247 -288 -3231 288
rect -3297 -300 -3231 -288
rect -3201 288 -3135 300
rect -3201 -288 -3185 288
rect -3151 -288 -3135 288
rect -3201 -300 -3135 -288
rect -3105 288 -3039 300
rect -3105 -288 -3089 288
rect -3055 -288 -3039 288
rect -3105 -300 -3039 -288
rect -3009 288 -2943 300
rect -3009 -288 -2993 288
rect -2959 -288 -2943 288
rect -3009 -300 -2943 -288
rect -2913 288 -2847 300
rect -2913 -288 -2897 288
rect -2863 -288 -2847 288
rect -2913 -300 -2847 -288
rect -2817 288 -2751 300
rect -2817 -288 -2801 288
rect -2767 -288 -2751 288
rect -2817 -300 -2751 -288
rect -2721 288 -2655 300
rect -2721 -288 -2705 288
rect -2671 -288 -2655 288
rect -2721 -300 -2655 -288
rect -2625 288 -2559 300
rect -2625 -288 -2609 288
rect -2575 -288 -2559 288
rect -2625 -300 -2559 -288
rect -2529 288 -2463 300
rect -2529 -288 -2513 288
rect -2479 -288 -2463 288
rect -2529 -300 -2463 -288
rect -2433 288 -2367 300
rect -2433 -288 -2417 288
rect -2383 -288 -2367 288
rect -2433 -300 -2367 -288
rect -2337 288 -2271 300
rect -2337 -288 -2321 288
rect -2287 -288 -2271 288
rect -2337 -300 -2271 -288
rect -2241 288 -2175 300
rect -2241 -288 -2225 288
rect -2191 -288 -2175 288
rect -2241 -300 -2175 -288
rect -2145 288 -2079 300
rect -2145 -288 -2129 288
rect -2095 -288 -2079 288
rect -2145 -300 -2079 -288
rect -2049 288 -1983 300
rect -2049 -288 -2033 288
rect -1999 -288 -1983 288
rect -2049 -300 -1983 -288
rect -1953 288 -1887 300
rect -1953 -288 -1937 288
rect -1903 -288 -1887 288
rect -1953 -300 -1887 -288
rect -1857 288 -1791 300
rect -1857 -288 -1841 288
rect -1807 -288 -1791 288
rect -1857 -300 -1791 -288
rect -1761 288 -1695 300
rect -1761 -288 -1745 288
rect -1711 -288 -1695 288
rect -1761 -300 -1695 -288
rect -1665 288 -1599 300
rect -1665 -288 -1649 288
rect -1615 -288 -1599 288
rect -1665 -300 -1599 -288
rect -1569 288 -1503 300
rect -1569 -288 -1553 288
rect -1519 -288 -1503 288
rect -1569 -300 -1503 -288
rect -1473 288 -1407 300
rect -1473 -288 -1457 288
rect -1423 -288 -1407 288
rect -1473 -300 -1407 -288
rect -1377 288 -1311 300
rect -1377 -288 -1361 288
rect -1327 -288 -1311 288
rect -1377 -300 -1311 -288
rect -1281 288 -1215 300
rect -1281 -288 -1265 288
rect -1231 -288 -1215 288
rect -1281 -300 -1215 -288
rect -1185 288 -1119 300
rect -1185 -288 -1169 288
rect -1135 -288 -1119 288
rect -1185 -300 -1119 -288
rect -1089 288 -1023 300
rect -1089 -288 -1073 288
rect -1039 -288 -1023 288
rect -1089 -300 -1023 -288
rect -993 288 -927 300
rect -993 -288 -977 288
rect -943 -288 -927 288
rect -993 -300 -927 -288
rect -897 288 -831 300
rect -897 -288 -881 288
rect -847 -288 -831 288
rect -897 -300 -831 -288
rect -801 288 -735 300
rect -801 -288 -785 288
rect -751 -288 -735 288
rect -801 -300 -735 -288
rect -705 288 -639 300
rect -705 -288 -689 288
rect -655 -288 -639 288
rect -705 -300 -639 -288
rect -609 288 -543 300
rect -609 -288 -593 288
rect -559 -288 -543 288
rect -609 -300 -543 -288
rect -513 288 -447 300
rect -513 -288 -497 288
rect -463 -288 -447 288
rect -513 -300 -447 -288
rect -417 288 -351 300
rect -417 -288 -401 288
rect -367 -288 -351 288
rect -417 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 417 300
rect 351 -288 367 288
rect 401 -288 417 288
rect 351 -300 417 -288
rect 447 288 513 300
rect 447 -288 463 288
rect 497 -288 513 288
rect 447 -300 513 -288
rect 543 288 609 300
rect 543 -288 559 288
rect 593 -288 609 288
rect 543 -300 609 -288
rect 639 288 705 300
rect 639 -288 655 288
rect 689 -288 705 288
rect 639 -300 705 -288
rect 735 288 801 300
rect 735 -288 751 288
rect 785 -288 801 288
rect 735 -300 801 -288
rect 831 288 897 300
rect 831 -288 847 288
rect 881 -288 897 288
rect 831 -300 897 -288
rect 927 288 993 300
rect 927 -288 943 288
rect 977 -288 993 288
rect 927 -300 993 -288
rect 1023 288 1089 300
rect 1023 -288 1039 288
rect 1073 -288 1089 288
rect 1023 -300 1089 -288
rect 1119 288 1185 300
rect 1119 -288 1135 288
rect 1169 -288 1185 288
rect 1119 -300 1185 -288
rect 1215 288 1281 300
rect 1215 -288 1231 288
rect 1265 -288 1281 288
rect 1215 -300 1281 -288
rect 1311 288 1377 300
rect 1311 -288 1327 288
rect 1361 -288 1377 288
rect 1311 -300 1377 -288
rect 1407 288 1473 300
rect 1407 -288 1423 288
rect 1457 -288 1473 288
rect 1407 -300 1473 -288
rect 1503 288 1569 300
rect 1503 -288 1519 288
rect 1553 -288 1569 288
rect 1503 -300 1569 -288
rect 1599 288 1665 300
rect 1599 -288 1615 288
rect 1649 -288 1665 288
rect 1599 -300 1665 -288
rect 1695 288 1761 300
rect 1695 -288 1711 288
rect 1745 -288 1761 288
rect 1695 -300 1761 -288
rect 1791 288 1857 300
rect 1791 -288 1807 288
rect 1841 -288 1857 288
rect 1791 -300 1857 -288
rect 1887 288 1953 300
rect 1887 -288 1903 288
rect 1937 -288 1953 288
rect 1887 -300 1953 -288
rect 1983 288 2049 300
rect 1983 -288 1999 288
rect 2033 -288 2049 288
rect 1983 -300 2049 -288
rect 2079 288 2145 300
rect 2079 -288 2095 288
rect 2129 -288 2145 288
rect 2079 -300 2145 -288
rect 2175 288 2241 300
rect 2175 -288 2191 288
rect 2225 -288 2241 288
rect 2175 -300 2241 -288
rect 2271 288 2337 300
rect 2271 -288 2287 288
rect 2321 -288 2337 288
rect 2271 -300 2337 -288
rect 2367 288 2433 300
rect 2367 -288 2383 288
rect 2417 -288 2433 288
rect 2367 -300 2433 -288
rect 2463 288 2529 300
rect 2463 -288 2479 288
rect 2513 -288 2529 288
rect 2463 -300 2529 -288
rect 2559 288 2625 300
rect 2559 -288 2575 288
rect 2609 -288 2625 288
rect 2559 -300 2625 -288
rect 2655 288 2721 300
rect 2655 -288 2671 288
rect 2705 -288 2721 288
rect 2655 -300 2721 -288
rect 2751 288 2817 300
rect 2751 -288 2767 288
rect 2801 -288 2817 288
rect 2751 -300 2817 -288
rect 2847 288 2913 300
rect 2847 -288 2863 288
rect 2897 -288 2913 288
rect 2847 -300 2913 -288
rect 2943 288 3009 300
rect 2943 -288 2959 288
rect 2993 -288 3009 288
rect 2943 -300 3009 -288
rect 3039 288 3105 300
rect 3039 -288 3055 288
rect 3089 -288 3105 288
rect 3039 -300 3105 -288
rect 3135 288 3201 300
rect 3135 -288 3151 288
rect 3185 -288 3201 288
rect 3135 -300 3201 -288
rect 3231 288 3297 300
rect 3231 -288 3247 288
rect 3281 -288 3297 288
rect 3231 -300 3297 -288
rect 3327 288 3393 300
rect 3327 -288 3343 288
rect 3377 -288 3393 288
rect 3327 -300 3393 -288
rect 3423 288 3489 300
rect 3423 -288 3439 288
rect 3473 -288 3489 288
rect 3423 -300 3489 -288
rect 3519 288 3585 300
rect 3519 -288 3535 288
rect 3569 -288 3585 288
rect 3519 -300 3585 -288
rect 3615 288 3681 300
rect 3615 -288 3631 288
rect 3665 -288 3681 288
rect 3615 -300 3681 -288
rect 3711 288 3777 300
rect 3711 -288 3727 288
rect 3761 -288 3777 288
rect 3711 -300 3777 -288
rect 3807 288 3873 300
rect 3807 -288 3823 288
rect 3857 -288 3873 288
rect 3807 -300 3873 -288
rect 3903 288 3969 300
rect 3903 -288 3919 288
rect 3953 -288 3969 288
rect 3903 -300 3969 -288
rect 3999 288 4065 300
rect 3999 -288 4015 288
rect 4049 -288 4065 288
rect 3999 -300 4065 -288
rect 4095 288 4161 300
rect 4095 -288 4111 288
rect 4145 -288 4161 288
rect 4095 -300 4161 -288
rect 4191 288 4257 300
rect 4191 -288 4207 288
rect 4241 -288 4257 288
rect 4191 -300 4257 -288
rect 4287 288 4349 300
rect 4287 -288 4303 288
rect 4337 -288 4349 288
rect 4287 -300 4349 -288
<< ndiffc >>
rect -4337 -288 -4303 288
rect -4241 -288 -4207 288
rect -4145 -288 -4111 288
rect -4049 -288 -4015 288
rect -3953 -288 -3919 288
rect -3857 -288 -3823 288
rect -3761 -288 -3727 288
rect -3665 -288 -3631 288
rect -3569 -288 -3535 288
rect -3473 -288 -3439 288
rect -3377 -288 -3343 288
rect -3281 -288 -3247 288
rect -3185 -288 -3151 288
rect -3089 -288 -3055 288
rect -2993 -288 -2959 288
rect -2897 -288 -2863 288
rect -2801 -288 -2767 288
rect -2705 -288 -2671 288
rect -2609 -288 -2575 288
rect -2513 -288 -2479 288
rect -2417 -288 -2383 288
rect -2321 -288 -2287 288
rect -2225 -288 -2191 288
rect -2129 -288 -2095 288
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
rect 2095 -288 2129 288
rect 2191 -288 2225 288
rect 2287 -288 2321 288
rect 2383 -288 2417 288
rect 2479 -288 2513 288
rect 2575 -288 2609 288
rect 2671 -288 2705 288
rect 2767 -288 2801 288
rect 2863 -288 2897 288
rect 2959 -288 2993 288
rect 3055 -288 3089 288
rect 3151 -288 3185 288
rect 3247 -288 3281 288
rect 3343 -288 3377 288
rect 3439 -288 3473 288
rect 3535 -288 3569 288
rect 3631 -288 3665 288
rect 3727 -288 3761 288
rect 3823 -288 3857 288
rect 3919 -288 3953 288
rect 4015 -288 4049 288
rect 4111 -288 4145 288
rect 4207 -288 4241 288
rect 4303 -288 4337 288
<< psubdiff >>
rect -4451 440 -4355 474
rect 4355 440 4451 474
rect -4451 378 -4417 440
rect 4417 378 4451 440
rect -4451 -440 -4417 -378
rect 4417 -440 4451 -378
rect -4451 -474 -4355 -440
rect 4355 -474 4451 -440
<< psubdiffcont >>
rect -4355 440 4355 474
rect -4451 -378 -4417 378
rect 4417 -378 4451 378
rect -4355 -474 4355 -440
<< poly >>
rect -4209 372 -4143 388
rect -4209 338 -4193 372
rect -4159 338 -4143 372
rect -4287 300 -4257 326
rect -4209 322 -4143 338
rect -4017 372 -3951 388
rect -4017 338 -4001 372
rect -3967 338 -3951 372
rect -4191 300 -4161 322
rect -4095 300 -4065 326
rect -4017 322 -3951 338
rect -3825 372 -3759 388
rect -3825 338 -3809 372
rect -3775 338 -3759 372
rect -3999 300 -3969 322
rect -3903 300 -3873 326
rect -3825 322 -3759 338
rect -3633 372 -3567 388
rect -3633 338 -3617 372
rect -3583 338 -3567 372
rect -3807 300 -3777 322
rect -3711 300 -3681 326
rect -3633 322 -3567 338
rect -3441 372 -3375 388
rect -3441 338 -3425 372
rect -3391 338 -3375 372
rect -3615 300 -3585 322
rect -3519 300 -3489 326
rect -3441 322 -3375 338
rect -3249 372 -3183 388
rect -3249 338 -3233 372
rect -3199 338 -3183 372
rect -3423 300 -3393 322
rect -3327 300 -3297 326
rect -3249 322 -3183 338
rect -3057 372 -2991 388
rect -3057 338 -3041 372
rect -3007 338 -2991 372
rect -3231 300 -3201 322
rect -3135 300 -3105 326
rect -3057 322 -2991 338
rect -2865 372 -2799 388
rect -2865 338 -2849 372
rect -2815 338 -2799 372
rect -3039 300 -3009 322
rect -2943 300 -2913 326
rect -2865 322 -2799 338
rect -2673 372 -2607 388
rect -2673 338 -2657 372
rect -2623 338 -2607 372
rect -2847 300 -2817 322
rect -2751 300 -2721 326
rect -2673 322 -2607 338
rect -2481 372 -2415 388
rect -2481 338 -2465 372
rect -2431 338 -2415 372
rect -2655 300 -2625 322
rect -2559 300 -2529 326
rect -2481 322 -2415 338
rect -2289 372 -2223 388
rect -2289 338 -2273 372
rect -2239 338 -2223 372
rect -2463 300 -2433 322
rect -2367 300 -2337 326
rect -2289 322 -2223 338
rect -2097 372 -2031 388
rect -2097 338 -2081 372
rect -2047 338 -2031 372
rect -2271 300 -2241 322
rect -2175 300 -2145 326
rect -2097 322 -2031 338
rect -1905 372 -1839 388
rect -1905 338 -1889 372
rect -1855 338 -1839 372
rect -2079 300 -2049 322
rect -1983 300 -1953 326
rect -1905 322 -1839 338
rect -1713 372 -1647 388
rect -1713 338 -1697 372
rect -1663 338 -1647 372
rect -1887 300 -1857 322
rect -1791 300 -1761 326
rect -1713 322 -1647 338
rect -1521 372 -1455 388
rect -1521 338 -1505 372
rect -1471 338 -1455 372
rect -1695 300 -1665 322
rect -1599 300 -1569 326
rect -1521 322 -1455 338
rect -1329 372 -1263 388
rect -1329 338 -1313 372
rect -1279 338 -1263 372
rect -1503 300 -1473 322
rect -1407 300 -1377 326
rect -1329 322 -1263 338
rect -1137 372 -1071 388
rect -1137 338 -1121 372
rect -1087 338 -1071 372
rect -1311 300 -1281 322
rect -1215 300 -1185 326
rect -1137 322 -1071 338
rect -945 372 -879 388
rect -945 338 -929 372
rect -895 338 -879 372
rect -1119 300 -1089 322
rect -1023 300 -993 326
rect -945 322 -879 338
rect -753 372 -687 388
rect -753 338 -737 372
rect -703 338 -687 372
rect -927 300 -897 322
rect -831 300 -801 326
rect -753 322 -687 338
rect -561 372 -495 388
rect -561 338 -545 372
rect -511 338 -495 372
rect -735 300 -705 322
rect -639 300 -609 326
rect -561 322 -495 338
rect -369 372 -303 388
rect -369 338 -353 372
rect -319 338 -303 372
rect -543 300 -513 322
rect -447 300 -417 326
rect -369 322 -303 338
rect -177 372 -111 388
rect -177 338 -161 372
rect -127 338 -111 372
rect -351 300 -321 322
rect -255 300 -225 326
rect -177 322 -111 338
rect 15 372 81 388
rect 15 338 31 372
rect 65 338 81 372
rect -159 300 -129 322
rect -63 300 -33 326
rect 15 322 81 338
rect 207 372 273 388
rect 207 338 223 372
rect 257 338 273 372
rect 33 300 63 322
rect 129 300 159 326
rect 207 322 273 338
rect 399 372 465 388
rect 399 338 415 372
rect 449 338 465 372
rect 225 300 255 322
rect 321 300 351 326
rect 399 322 465 338
rect 591 372 657 388
rect 591 338 607 372
rect 641 338 657 372
rect 417 300 447 322
rect 513 300 543 326
rect 591 322 657 338
rect 783 372 849 388
rect 783 338 799 372
rect 833 338 849 372
rect 609 300 639 322
rect 705 300 735 326
rect 783 322 849 338
rect 975 372 1041 388
rect 975 338 991 372
rect 1025 338 1041 372
rect 801 300 831 322
rect 897 300 927 326
rect 975 322 1041 338
rect 1167 372 1233 388
rect 1167 338 1183 372
rect 1217 338 1233 372
rect 993 300 1023 322
rect 1089 300 1119 326
rect 1167 322 1233 338
rect 1359 372 1425 388
rect 1359 338 1375 372
rect 1409 338 1425 372
rect 1185 300 1215 322
rect 1281 300 1311 326
rect 1359 322 1425 338
rect 1551 372 1617 388
rect 1551 338 1567 372
rect 1601 338 1617 372
rect 1377 300 1407 322
rect 1473 300 1503 326
rect 1551 322 1617 338
rect 1743 372 1809 388
rect 1743 338 1759 372
rect 1793 338 1809 372
rect 1569 300 1599 322
rect 1665 300 1695 326
rect 1743 322 1809 338
rect 1935 372 2001 388
rect 1935 338 1951 372
rect 1985 338 2001 372
rect 1761 300 1791 322
rect 1857 300 1887 326
rect 1935 322 2001 338
rect 2127 372 2193 388
rect 2127 338 2143 372
rect 2177 338 2193 372
rect 1953 300 1983 322
rect 2049 300 2079 326
rect 2127 322 2193 338
rect 2319 372 2385 388
rect 2319 338 2335 372
rect 2369 338 2385 372
rect 2145 300 2175 322
rect 2241 300 2271 326
rect 2319 322 2385 338
rect 2511 372 2577 388
rect 2511 338 2527 372
rect 2561 338 2577 372
rect 2337 300 2367 322
rect 2433 300 2463 326
rect 2511 322 2577 338
rect 2703 372 2769 388
rect 2703 338 2719 372
rect 2753 338 2769 372
rect 2529 300 2559 322
rect 2625 300 2655 326
rect 2703 322 2769 338
rect 2895 372 2961 388
rect 2895 338 2911 372
rect 2945 338 2961 372
rect 2721 300 2751 322
rect 2817 300 2847 326
rect 2895 322 2961 338
rect 3087 372 3153 388
rect 3087 338 3103 372
rect 3137 338 3153 372
rect 2913 300 2943 322
rect 3009 300 3039 326
rect 3087 322 3153 338
rect 3279 372 3345 388
rect 3279 338 3295 372
rect 3329 338 3345 372
rect 3105 300 3135 322
rect 3201 300 3231 326
rect 3279 322 3345 338
rect 3471 372 3537 388
rect 3471 338 3487 372
rect 3521 338 3537 372
rect 3297 300 3327 322
rect 3393 300 3423 326
rect 3471 322 3537 338
rect 3663 372 3729 388
rect 3663 338 3679 372
rect 3713 338 3729 372
rect 3489 300 3519 322
rect 3585 300 3615 326
rect 3663 322 3729 338
rect 3855 372 3921 388
rect 3855 338 3871 372
rect 3905 338 3921 372
rect 3681 300 3711 322
rect 3777 300 3807 326
rect 3855 322 3921 338
rect 4047 372 4113 388
rect 4047 338 4063 372
rect 4097 338 4113 372
rect 3873 300 3903 322
rect 3969 300 3999 326
rect 4047 322 4113 338
rect 4239 372 4305 388
rect 4239 338 4255 372
rect 4289 338 4305 372
rect 4065 300 4095 322
rect 4161 300 4191 326
rect 4239 322 4305 338
rect 4257 300 4287 322
rect -4287 -322 -4257 -300
rect -4305 -338 -4239 -322
rect -4191 -326 -4161 -300
rect -4095 -322 -4065 -300
rect -4305 -372 -4289 -338
rect -4255 -372 -4239 -338
rect -4305 -388 -4239 -372
rect -4113 -338 -4047 -322
rect -3999 -326 -3969 -300
rect -3903 -322 -3873 -300
rect -4113 -372 -4097 -338
rect -4063 -372 -4047 -338
rect -4113 -388 -4047 -372
rect -3921 -338 -3855 -322
rect -3807 -326 -3777 -300
rect -3711 -322 -3681 -300
rect -3921 -372 -3905 -338
rect -3871 -372 -3855 -338
rect -3921 -388 -3855 -372
rect -3729 -338 -3663 -322
rect -3615 -326 -3585 -300
rect -3519 -322 -3489 -300
rect -3729 -372 -3713 -338
rect -3679 -372 -3663 -338
rect -3729 -388 -3663 -372
rect -3537 -338 -3471 -322
rect -3423 -326 -3393 -300
rect -3327 -322 -3297 -300
rect -3537 -372 -3521 -338
rect -3487 -372 -3471 -338
rect -3537 -388 -3471 -372
rect -3345 -338 -3279 -322
rect -3231 -326 -3201 -300
rect -3135 -322 -3105 -300
rect -3345 -372 -3329 -338
rect -3295 -372 -3279 -338
rect -3345 -388 -3279 -372
rect -3153 -338 -3087 -322
rect -3039 -326 -3009 -300
rect -2943 -322 -2913 -300
rect -3153 -372 -3137 -338
rect -3103 -372 -3087 -338
rect -3153 -388 -3087 -372
rect -2961 -338 -2895 -322
rect -2847 -326 -2817 -300
rect -2751 -322 -2721 -300
rect -2961 -372 -2945 -338
rect -2911 -372 -2895 -338
rect -2961 -388 -2895 -372
rect -2769 -338 -2703 -322
rect -2655 -326 -2625 -300
rect -2559 -322 -2529 -300
rect -2769 -372 -2753 -338
rect -2719 -372 -2703 -338
rect -2769 -388 -2703 -372
rect -2577 -338 -2511 -322
rect -2463 -326 -2433 -300
rect -2367 -322 -2337 -300
rect -2577 -372 -2561 -338
rect -2527 -372 -2511 -338
rect -2577 -388 -2511 -372
rect -2385 -338 -2319 -322
rect -2271 -326 -2241 -300
rect -2175 -322 -2145 -300
rect -2385 -372 -2369 -338
rect -2335 -372 -2319 -338
rect -2385 -388 -2319 -372
rect -2193 -338 -2127 -322
rect -2079 -326 -2049 -300
rect -1983 -322 -1953 -300
rect -2193 -372 -2177 -338
rect -2143 -372 -2127 -338
rect -2193 -388 -2127 -372
rect -2001 -338 -1935 -322
rect -1887 -326 -1857 -300
rect -1791 -322 -1761 -300
rect -2001 -372 -1985 -338
rect -1951 -372 -1935 -338
rect -2001 -388 -1935 -372
rect -1809 -338 -1743 -322
rect -1695 -326 -1665 -300
rect -1599 -322 -1569 -300
rect -1809 -372 -1793 -338
rect -1759 -372 -1743 -338
rect -1809 -388 -1743 -372
rect -1617 -338 -1551 -322
rect -1503 -326 -1473 -300
rect -1407 -322 -1377 -300
rect -1617 -372 -1601 -338
rect -1567 -372 -1551 -338
rect -1617 -388 -1551 -372
rect -1425 -338 -1359 -322
rect -1311 -326 -1281 -300
rect -1215 -322 -1185 -300
rect -1425 -372 -1409 -338
rect -1375 -372 -1359 -338
rect -1425 -388 -1359 -372
rect -1233 -338 -1167 -322
rect -1119 -326 -1089 -300
rect -1023 -322 -993 -300
rect -1233 -372 -1217 -338
rect -1183 -372 -1167 -338
rect -1233 -388 -1167 -372
rect -1041 -338 -975 -322
rect -927 -326 -897 -300
rect -831 -322 -801 -300
rect -1041 -372 -1025 -338
rect -991 -372 -975 -338
rect -1041 -388 -975 -372
rect -849 -338 -783 -322
rect -735 -326 -705 -300
rect -639 -322 -609 -300
rect -849 -372 -833 -338
rect -799 -372 -783 -338
rect -849 -388 -783 -372
rect -657 -338 -591 -322
rect -543 -326 -513 -300
rect -447 -322 -417 -300
rect -657 -372 -641 -338
rect -607 -372 -591 -338
rect -657 -388 -591 -372
rect -465 -338 -399 -322
rect -351 -326 -321 -300
rect -255 -322 -225 -300
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -465 -388 -399 -372
rect -273 -338 -207 -322
rect -159 -326 -129 -300
rect -63 -322 -33 -300
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -273 -388 -207 -372
rect -81 -338 -15 -322
rect 33 -326 63 -300
rect 129 -322 159 -300
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect -81 -388 -15 -372
rect 111 -338 177 -322
rect 225 -326 255 -300
rect 321 -322 351 -300
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 111 -388 177 -372
rect 303 -338 369 -322
rect 417 -326 447 -300
rect 513 -322 543 -300
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 303 -388 369 -372
rect 495 -338 561 -322
rect 609 -326 639 -300
rect 705 -322 735 -300
rect 495 -372 511 -338
rect 545 -372 561 -338
rect 495 -388 561 -372
rect 687 -338 753 -322
rect 801 -326 831 -300
rect 897 -322 927 -300
rect 687 -372 703 -338
rect 737 -372 753 -338
rect 687 -388 753 -372
rect 879 -338 945 -322
rect 993 -326 1023 -300
rect 1089 -322 1119 -300
rect 879 -372 895 -338
rect 929 -372 945 -338
rect 879 -388 945 -372
rect 1071 -338 1137 -322
rect 1185 -326 1215 -300
rect 1281 -322 1311 -300
rect 1071 -372 1087 -338
rect 1121 -372 1137 -338
rect 1071 -388 1137 -372
rect 1263 -338 1329 -322
rect 1377 -326 1407 -300
rect 1473 -322 1503 -300
rect 1263 -372 1279 -338
rect 1313 -372 1329 -338
rect 1263 -388 1329 -372
rect 1455 -338 1521 -322
rect 1569 -326 1599 -300
rect 1665 -322 1695 -300
rect 1455 -372 1471 -338
rect 1505 -372 1521 -338
rect 1455 -388 1521 -372
rect 1647 -338 1713 -322
rect 1761 -326 1791 -300
rect 1857 -322 1887 -300
rect 1647 -372 1663 -338
rect 1697 -372 1713 -338
rect 1647 -388 1713 -372
rect 1839 -338 1905 -322
rect 1953 -326 1983 -300
rect 2049 -322 2079 -300
rect 1839 -372 1855 -338
rect 1889 -372 1905 -338
rect 1839 -388 1905 -372
rect 2031 -338 2097 -322
rect 2145 -326 2175 -300
rect 2241 -322 2271 -300
rect 2031 -372 2047 -338
rect 2081 -372 2097 -338
rect 2031 -388 2097 -372
rect 2223 -338 2289 -322
rect 2337 -326 2367 -300
rect 2433 -322 2463 -300
rect 2223 -372 2239 -338
rect 2273 -372 2289 -338
rect 2223 -388 2289 -372
rect 2415 -338 2481 -322
rect 2529 -326 2559 -300
rect 2625 -322 2655 -300
rect 2415 -372 2431 -338
rect 2465 -372 2481 -338
rect 2415 -388 2481 -372
rect 2607 -338 2673 -322
rect 2721 -326 2751 -300
rect 2817 -322 2847 -300
rect 2607 -372 2623 -338
rect 2657 -372 2673 -338
rect 2607 -388 2673 -372
rect 2799 -338 2865 -322
rect 2913 -326 2943 -300
rect 3009 -322 3039 -300
rect 2799 -372 2815 -338
rect 2849 -372 2865 -338
rect 2799 -388 2865 -372
rect 2991 -338 3057 -322
rect 3105 -326 3135 -300
rect 3201 -322 3231 -300
rect 2991 -372 3007 -338
rect 3041 -372 3057 -338
rect 2991 -388 3057 -372
rect 3183 -338 3249 -322
rect 3297 -326 3327 -300
rect 3393 -322 3423 -300
rect 3183 -372 3199 -338
rect 3233 -372 3249 -338
rect 3183 -388 3249 -372
rect 3375 -338 3441 -322
rect 3489 -326 3519 -300
rect 3585 -322 3615 -300
rect 3375 -372 3391 -338
rect 3425 -372 3441 -338
rect 3375 -388 3441 -372
rect 3567 -338 3633 -322
rect 3681 -326 3711 -300
rect 3777 -322 3807 -300
rect 3567 -372 3583 -338
rect 3617 -372 3633 -338
rect 3567 -388 3633 -372
rect 3759 -338 3825 -322
rect 3873 -326 3903 -300
rect 3969 -322 3999 -300
rect 3759 -372 3775 -338
rect 3809 -372 3825 -338
rect 3759 -388 3825 -372
rect 3951 -338 4017 -322
rect 4065 -326 4095 -300
rect 4161 -322 4191 -300
rect 3951 -372 3967 -338
rect 4001 -372 4017 -338
rect 3951 -388 4017 -372
rect 4143 -338 4209 -322
rect 4257 -326 4287 -300
rect 4143 -372 4159 -338
rect 4193 -372 4209 -338
rect 4143 -388 4209 -372
<< polycont >>
rect -4193 338 -4159 372
rect -4001 338 -3967 372
rect -3809 338 -3775 372
rect -3617 338 -3583 372
rect -3425 338 -3391 372
rect -3233 338 -3199 372
rect -3041 338 -3007 372
rect -2849 338 -2815 372
rect -2657 338 -2623 372
rect -2465 338 -2431 372
rect -2273 338 -2239 372
rect -2081 338 -2047 372
rect -1889 338 -1855 372
rect -1697 338 -1663 372
rect -1505 338 -1471 372
rect -1313 338 -1279 372
rect -1121 338 -1087 372
rect -929 338 -895 372
rect -737 338 -703 372
rect -545 338 -511 372
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect 607 338 641 372
rect 799 338 833 372
rect 991 338 1025 372
rect 1183 338 1217 372
rect 1375 338 1409 372
rect 1567 338 1601 372
rect 1759 338 1793 372
rect 1951 338 1985 372
rect 2143 338 2177 372
rect 2335 338 2369 372
rect 2527 338 2561 372
rect 2719 338 2753 372
rect 2911 338 2945 372
rect 3103 338 3137 372
rect 3295 338 3329 372
rect 3487 338 3521 372
rect 3679 338 3713 372
rect 3871 338 3905 372
rect 4063 338 4097 372
rect 4255 338 4289 372
rect -4289 -372 -4255 -338
rect -4097 -372 -4063 -338
rect -3905 -372 -3871 -338
rect -3713 -372 -3679 -338
rect -3521 -372 -3487 -338
rect -3329 -372 -3295 -338
rect -3137 -372 -3103 -338
rect -2945 -372 -2911 -338
rect -2753 -372 -2719 -338
rect -2561 -372 -2527 -338
rect -2369 -372 -2335 -338
rect -2177 -372 -2143 -338
rect -1985 -372 -1951 -338
rect -1793 -372 -1759 -338
rect -1601 -372 -1567 -338
rect -1409 -372 -1375 -338
rect -1217 -372 -1183 -338
rect -1025 -372 -991 -338
rect -833 -372 -799 -338
rect -641 -372 -607 -338
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
rect 511 -372 545 -338
rect 703 -372 737 -338
rect 895 -372 929 -338
rect 1087 -372 1121 -338
rect 1279 -372 1313 -338
rect 1471 -372 1505 -338
rect 1663 -372 1697 -338
rect 1855 -372 1889 -338
rect 2047 -372 2081 -338
rect 2239 -372 2273 -338
rect 2431 -372 2465 -338
rect 2623 -372 2657 -338
rect 2815 -372 2849 -338
rect 3007 -372 3041 -338
rect 3199 -372 3233 -338
rect 3391 -372 3425 -338
rect 3583 -372 3617 -338
rect 3775 -372 3809 -338
rect 3967 -372 4001 -338
rect 4159 -372 4193 -338
<< locali >>
rect -4451 440 -4355 474
rect 4355 440 4451 474
rect -4451 378 -4417 440
rect 4417 378 4451 440
rect -4209 338 -4193 372
rect -4159 338 -4143 372
rect -4017 338 -4001 372
rect -3967 338 -3951 372
rect -3825 338 -3809 372
rect -3775 338 -3759 372
rect -3633 338 -3617 372
rect -3583 338 -3567 372
rect -3441 338 -3425 372
rect -3391 338 -3375 372
rect -3249 338 -3233 372
rect -3199 338 -3183 372
rect -3057 338 -3041 372
rect -3007 338 -2991 372
rect -2865 338 -2849 372
rect -2815 338 -2799 372
rect -2673 338 -2657 372
rect -2623 338 -2607 372
rect -2481 338 -2465 372
rect -2431 338 -2415 372
rect -2289 338 -2273 372
rect -2239 338 -2223 372
rect -2097 338 -2081 372
rect -2047 338 -2031 372
rect -1905 338 -1889 372
rect -1855 338 -1839 372
rect -1713 338 -1697 372
rect -1663 338 -1647 372
rect -1521 338 -1505 372
rect -1471 338 -1455 372
rect -1329 338 -1313 372
rect -1279 338 -1263 372
rect -1137 338 -1121 372
rect -1087 338 -1071 372
rect -945 338 -929 372
rect -895 338 -879 372
rect -753 338 -737 372
rect -703 338 -687 372
rect -561 338 -545 372
rect -511 338 -495 372
rect -369 338 -353 372
rect -319 338 -303 372
rect -177 338 -161 372
rect -127 338 -111 372
rect 15 338 31 372
rect 65 338 81 372
rect 207 338 223 372
rect 257 338 273 372
rect 399 338 415 372
rect 449 338 465 372
rect 591 338 607 372
rect 641 338 657 372
rect 783 338 799 372
rect 833 338 849 372
rect 975 338 991 372
rect 1025 338 1041 372
rect 1167 338 1183 372
rect 1217 338 1233 372
rect 1359 338 1375 372
rect 1409 338 1425 372
rect 1551 338 1567 372
rect 1601 338 1617 372
rect 1743 338 1759 372
rect 1793 338 1809 372
rect 1935 338 1951 372
rect 1985 338 2001 372
rect 2127 338 2143 372
rect 2177 338 2193 372
rect 2319 338 2335 372
rect 2369 338 2385 372
rect 2511 338 2527 372
rect 2561 338 2577 372
rect 2703 338 2719 372
rect 2753 338 2769 372
rect 2895 338 2911 372
rect 2945 338 2961 372
rect 3087 338 3103 372
rect 3137 338 3153 372
rect 3279 338 3295 372
rect 3329 338 3345 372
rect 3471 338 3487 372
rect 3521 338 3537 372
rect 3663 338 3679 372
rect 3713 338 3729 372
rect 3855 338 3871 372
rect 3905 338 3921 372
rect 4047 338 4063 372
rect 4097 338 4113 372
rect 4239 338 4255 372
rect 4289 338 4305 372
rect -4337 288 -4303 304
rect -4337 -304 -4303 -288
rect -4241 288 -4207 304
rect -4241 -304 -4207 -288
rect -4145 288 -4111 304
rect -4145 -304 -4111 -288
rect -4049 288 -4015 304
rect -4049 -304 -4015 -288
rect -3953 288 -3919 304
rect -3953 -304 -3919 -288
rect -3857 288 -3823 304
rect -3857 -304 -3823 -288
rect -3761 288 -3727 304
rect -3761 -304 -3727 -288
rect -3665 288 -3631 304
rect -3665 -304 -3631 -288
rect -3569 288 -3535 304
rect -3569 -304 -3535 -288
rect -3473 288 -3439 304
rect -3473 -304 -3439 -288
rect -3377 288 -3343 304
rect -3377 -304 -3343 -288
rect -3281 288 -3247 304
rect -3281 -304 -3247 -288
rect -3185 288 -3151 304
rect -3185 -304 -3151 -288
rect -3089 288 -3055 304
rect -3089 -304 -3055 -288
rect -2993 288 -2959 304
rect -2993 -304 -2959 -288
rect -2897 288 -2863 304
rect -2897 -304 -2863 -288
rect -2801 288 -2767 304
rect -2801 -304 -2767 -288
rect -2705 288 -2671 304
rect -2705 -304 -2671 -288
rect -2609 288 -2575 304
rect -2609 -304 -2575 -288
rect -2513 288 -2479 304
rect -2513 -304 -2479 -288
rect -2417 288 -2383 304
rect -2417 -304 -2383 -288
rect -2321 288 -2287 304
rect -2321 -304 -2287 -288
rect -2225 288 -2191 304
rect -2225 -304 -2191 -288
rect -2129 288 -2095 304
rect -2129 -304 -2095 -288
rect -2033 288 -1999 304
rect -2033 -304 -1999 -288
rect -1937 288 -1903 304
rect -1937 -304 -1903 -288
rect -1841 288 -1807 304
rect -1841 -304 -1807 -288
rect -1745 288 -1711 304
rect -1745 -304 -1711 -288
rect -1649 288 -1615 304
rect -1649 -304 -1615 -288
rect -1553 288 -1519 304
rect -1553 -304 -1519 -288
rect -1457 288 -1423 304
rect -1457 -304 -1423 -288
rect -1361 288 -1327 304
rect -1361 -304 -1327 -288
rect -1265 288 -1231 304
rect -1265 -304 -1231 -288
rect -1169 288 -1135 304
rect -1169 -304 -1135 -288
rect -1073 288 -1039 304
rect -1073 -304 -1039 -288
rect -977 288 -943 304
rect -977 -304 -943 -288
rect -881 288 -847 304
rect -881 -304 -847 -288
rect -785 288 -751 304
rect -785 -304 -751 -288
rect -689 288 -655 304
rect -689 -304 -655 -288
rect -593 288 -559 304
rect -593 -304 -559 -288
rect -497 288 -463 304
rect -497 -304 -463 -288
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect 463 288 497 304
rect 463 -304 497 -288
rect 559 288 593 304
rect 559 -304 593 -288
rect 655 288 689 304
rect 655 -304 689 -288
rect 751 288 785 304
rect 751 -304 785 -288
rect 847 288 881 304
rect 847 -304 881 -288
rect 943 288 977 304
rect 943 -304 977 -288
rect 1039 288 1073 304
rect 1039 -304 1073 -288
rect 1135 288 1169 304
rect 1135 -304 1169 -288
rect 1231 288 1265 304
rect 1231 -304 1265 -288
rect 1327 288 1361 304
rect 1327 -304 1361 -288
rect 1423 288 1457 304
rect 1423 -304 1457 -288
rect 1519 288 1553 304
rect 1519 -304 1553 -288
rect 1615 288 1649 304
rect 1615 -304 1649 -288
rect 1711 288 1745 304
rect 1711 -304 1745 -288
rect 1807 288 1841 304
rect 1807 -304 1841 -288
rect 1903 288 1937 304
rect 1903 -304 1937 -288
rect 1999 288 2033 304
rect 1999 -304 2033 -288
rect 2095 288 2129 304
rect 2095 -304 2129 -288
rect 2191 288 2225 304
rect 2191 -304 2225 -288
rect 2287 288 2321 304
rect 2287 -304 2321 -288
rect 2383 288 2417 304
rect 2383 -304 2417 -288
rect 2479 288 2513 304
rect 2479 -304 2513 -288
rect 2575 288 2609 304
rect 2575 -304 2609 -288
rect 2671 288 2705 304
rect 2671 -304 2705 -288
rect 2767 288 2801 304
rect 2767 -304 2801 -288
rect 2863 288 2897 304
rect 2863 -304 2897 -288
rect 2959 288 2993 304
rect 2959 -304 2993 -288
rect 3055 288 3089 304
rect 3055 -304 3089 -288
rect 3151 288 3185 304
rect 3151 -304 3185 -288
rect 3247 288 3281 304
rect 3247 -304 3281 -288
rect 3343 288 3377 304
rect 3343 -304 3377 -288
rect 3439 288 3473 304
rect 3439 -304 3473 -288
rect 3535 288 3569 304
rect 3535 -304 3569 -288
rect 3631 288 3665 304
rect 3631 -304 3665 -288
rect 3727 288 3761 304
rect 3727 -304 3761 -288
rect 3823 288 3857 304
rect 3823 -304 3857 -288
rect 3919 288 3953 304
rect 3919 -304 3953 -288
rect 4015 288 4049 304
rect 4015 -304 4049 -288
rect 4111 288 4145 304
rect 4111 -304 4145 -288
rect 4207 288 4241 304
rect 4207 -304 4241 -288
rect 4303 288 4337 304
rect 4303 -304 4337 -288
rect -4305 -372 -4289 -338
rect -4255 -372 -4239 -338
rect -4113 -372 -4097 -338
rect -4063 -372 -4047 -338
rect -3921 -372 -3905 -338
rect -3871 -372 -3855 -338
rect -3729 -372 -3713 -338
rect -3679 -372 -3663 -338
rect -3537 -372 -3521 -338
rect -3487 -372 -3471 -338
rect -3345 -372 -3329 -338
rect -3295 -372 -3279 -338
rect -3153 -372 -3137 -338
rect -3103 -372 -3087 -338
rect -2961 -372 -2945 -338
rect -2911 -372 -2895 -338
rect -2769 -372 -2753 -338
rect -2719 -372 -2703 -338
rect -2577 -372 -2561 -338
rect -2527 -372 -2511 -338
rect -2385 -372 -2369 -338
rect -2335 -372 -2319 -338
rect -2193 -372 -2177 -338
rect -2143 -372 -2127 -338
rect -2001 -372 -1985 -338
rect -1951 -372 -1935 -338
rect -1809 -372 -1793 -338
rect -1759 -372 -1743 -338
rect -1617 -372 -1601 -338
rect -1567 -372 -1551 -338
rect -1425 -372 -1409 -338
rect -1375 -372 -1359 -338
rect -1233 -372 -1217 -338
rect -1183 -372 -1167 -338
rect -1041 -372 -1025 -338
rect -991 -372 -975 -338
rect -849 -372 -833 -338
rect -799 -372 -783 -338
rect -657 -372 -641 -338
rect -607 -372 -591 -338
rect -465 -372 -449 -338
rect -415 -372 -399 -338
rect -273 -372 -257 -338
rect -223 -372 -207 -338
rect -81 -372 -65 -338
rect -31 -372 -15 -338
rect 111 -372 127 -338
rect 161 -372 177 -338
rect 303 -372 319 -338
rect 353 -372 369 -338
rect 495 -372 511 -338
rect 545 -372 561 -338
rect 687 -372 703 -338
rect 737 -372 753 -338
rect 879 -372 895 -338
rect 929 -372 945 -338
rect 1071 -372 1087 -338
rect 1121 -372 1137 -338
rect 1263 -372 1279 -338
rect 1313 -372 1329 -338
rect 1455 -372 1471 -338
rect 1505 -372 1521 -338
rect 1647 -372 1663 -338
rect 1697 -372 1713 -338
rect 1839 -372 1855 -338
rect 1889 -372 1905 -338
rect 2031 -372 2047 -338
rect 2081 -372 2097 -338
rect 2223 -372 2239 -338
rect 2273 -372 2289 -338
rect 2415 -372 2431 -338
rect 2465 -372 2481 -338
rect 2607 -372 2623 -338
rect 2657 -372 2673 -338
rect 2799 -372 2815 -338
rect 2849 -372 2865 -338
rect 2991 -372 3007 -338
rect 3041 -372 3057 -338
rect 3183 -372 3199 -338
rect 3233 -372 3249 -338
rect 3375 -372 3391 -338
rect 3425 -372 3441 -338
rect 3567 -372 3583 -338
rect 3617 -372 3633 -338
rect 3759 -372 3775 -338
rect 3809 -372 3825 -338
rect 3951 -372 3967 -338
rect 4001 -372 4017 -338
rect 4143 -372 4159 -338
rect 4193 -372 4209 -338
rect -4451 -440 -4417 -378
rect 4417 -440 4451 -378
rect -4451 -474 -4355 -440
rect 4355 -474 4451 -440
<< viali >>
rect -4193 338 -4159 372
rect -4001 338 -3967 372
rect -3809 338 -3775 372
rect -3617 338 -3583 372
rect -3425 338 -3391 372
rect -3233 338 -3199 372
rect -3041 338 -3007 372
rect -2849 338 -2815 372
rect -2657 338 -2623 372
rect -2465 338 -2431 372
rect -2273 338 -2239 372
rect -2081 338 -2047 372
rect -1889 338 -1855 372
rect -1697 338 -1663 372
rect -1505 338 -1471 372
rect -1313 338 -1279 372
rect -1121 338 -1087 372
rect -929 338 -895 372
rect -737 338 -703 372
rect -545 338 -511 372
rect -353 338 -319 372
rect -161 338 -127 372
rect 31 338 65 372
rect 223 338 257 372
rect 415 338 449 372
rect 607 338 641 372
rect 799 338 833 372
rect 991 338 1025 372
rect 1183 338 1217 372
rect 1375 338 1409 372
rect 1567 338 1601 372
rect 1759 338 1793 372
rect 1951 338 1985 372
rect 2143 338 2177 372
rect 2335 338 2369 372
rect 2527 338 2561 372
rect 2719 338 2753 372
rect 2911 338 2945 372
rect 3103 338 3137 372
rect 3295 338 3329 372
rect 3487 338 3521 372
rect 3679 338 3713 372
rect 3871 338 3905 372
rect 4063 338 4097 372
rect 4255 338 4289 372
rect -4337 -288 -4303 288
rect -4241 -288 -4207 288
rect -4145 -288 -4111 288
rect -4049 -288 -4015 288
rect -3953 -288 -3919 288
rect -3857 -288 -3823 288
rect -3761 -288 -3727 288
rect -3665 -288 -3631 288
rect -3569 -288 -3535 288
rect -3473 -288 -3439 288
rect -3377 -288 -3343 288
rect -3281 -288 -3247 288
rect -3185 -288 -3151 288
rect -3089 -288 -3055 288
rect -2993 -288 -2959 288
rect -2897 -288 -2863 288
rect -2801 -288 -2767 288
rect -2705 -288 -2671 288
rect -2609 -288 -2575 288
rect -2513 -288 -2479 288
rect -2417 -288 -2383 288
rect -2321 -288 -2287 288
rect -2225 -288 -2191 288
rect -2129 -288 -2095 288
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
rect 2095 -288 2129 288
rect 2191 -288 2225 288
rect 2287 -288 2321 288
rect 2383 -288 2417 288
rect 2479 -288 2513 288
rect 2575 -288 2609 288
rect 2671 -288 2705 288
rect 2767 -288 2801 288
rect 2863 -288 2897 288
rect 2959 -288 2993 288
rect 3055 -288 3089 288
rect 3151 -288 3185 288
rect 3247 -288 3281 288
rect 3343 -288 3377 288
rect 3439 -288 3473 288
rect 3535 -288 3569 288
rect 3631 -288 3665 288
rect 3727 -288 3761 288
rect 3823 -288 3857 288
rect 3919 -288 3953 288
rect 4015 -288 4049 288
rect 4111 -288 4145 288
rect 4207 -288 4241 288
rect 4303 -288 4337 288
rect -4289 -372 -4255 -338
rect -4097 -372 -4063 -338
rect -3905 -372 -3871 -338
rect -3713 -372 -3679 -338
rect -3521 -372 -3487 -338
rect -3329 -372 -3295 -338
rect -3137 -372 -3103 -338
rect -2945 -372 -2911 -338
rect -2753 -372 -2719 -338
rect -2561 -372 -2527 -338
rect -2369 -372 -2335 -338
rect -2177 -372 -2143 -338
rect -1985 -372 -1951 -338
rect -1793 -372 -1759 -338
rect -1601 -372 -1567 -338
rect -1409 -372 -1375 -338
rect -1217 -372 -1183 -338
rect -1025 -372 -991 -338
rect -833 -372 -799 -338
rect -641 -372 -607 -338
rect -449 -372 -415 -338
rect -257 -372 -223 -338
rect -65 -372 -31 -338
rect 127 -372 161 -338
rect 319 -372 353 -338
rect 511 -372 545 -338
rect 703 -372 737 -338
rect 895 -372 929 -338
rect 1087 -372 1121 -338
rect 1279 -372 1313 -338
rect 1471 -372 1505 -338
rect 1663 -372 1697 -338
rect 1855 -372 1889 -338
rect 2047 -372 2081 -338
rect 2239 -372 2273 -338
rect 2431 -372 2465 -338
rect 2623 -372 2657 -338
rect 2815 -372 2849 -338
rect 3007 -372 3041 -338
rect 3199 -372 3233 -338
rect 3391 -372 3425 -338
rect 3583 -372 3617 -338
rect 3775 -372 3809 -338
rect 3967 -372 4001 -338
rect 4159 -372 4193 -338
<< metal1 >>
rect -4205 372 -4147 378
rect -4205 338 -4193 372
rect -4159 338 -4147 372
rect -4205 332 -4147 338
rect -4013 372 -3955 378
rect -4013 338 -4001 372
rect -3967 338 -3955 372
rect -4013 332 -3955 338
rect -3821 372 -3763 378
rect -3821 338 -3809 372
rect -3775 338 -3763 372
rect -3821 332 -3763 338
rect -3629 372 -3571 378
rect -3629 338 -3617 372
rect -3583 338 -3571 372
rect -3629 332 -3571 338
rect -3437 372 -3379 378
rect -3437 338 -3425 372
rect -3391 338 -3379 372
rect -3437 332 -3379 338
rect -3245 372 -3187 378
rect -3245 338 -3233 372
rect -3199 338 -3187 372
rect -3245 332 -3187 338
rect -3053 372 -2995 378
rect -3053 338 -3041 372
rect -3007 338 -2995 372
rect -3053 332 -2995 338
rect -2861 372 -2803 378
rect -2861 338 -2849 372
rect -2815 338 -2803 372
rect -2861 332 -2803 338
rect -2669 372 -2611 378
rect -2669 338 -2657 372
rect -2623 338 -2611 372
rect -2669 332 -2611 338
rect -2477 372 -2419 378
rect -2477 338 -2465 372
rect -2431 338 -2419 372
rect -2477 332 -2419 338
rect -2285 372 -2227 378
rect -2285 338 -2273 372
rect -2239 338 -2227 372
rect -2285 332 -2227 338
rect -2093 372 -2035 378
rect -2093 338 -2081 372
rect -2047 338 -2035 372
rect -2093 332 -2035 338
rect -1901 372 -1843 378
rect -1901 338 -1889 372
rect -1855 338 -1843 372
rect -1901 332 -1843 338
rect -1709 372 -1651 378
rect -1709 338 -1697 372
rect -1663 338 -1651 372
rect -1709 332 -1651 338
rect -1517 372 -1459 378
rect -1517 338 -1505 372
rect -1471 338 -1459 372
rect -1517 332 -1459 338
rect -1325 372 -1267 378
rect -1325 338 -1313 372
rect -1279 338 -1267 372
rect -1325 332 -1267 338
rect -1133 372 -1075 378
rect -1133 338 -1121 372
rect -1087 338 -1075 372
rect -1133 332 -1075 338
rect -941 372 -883 378
rect -941 338 -929 372
rect -895 338 -883 372
rect -941 332 -883 338
rect -749 372 -691 378
rect -749 338 -737 372
rect -703 338 -691 372
rect -749 332 -691 338
rect -557 372 -499 378
rect -557 338 -545 372
rect -511 338 -499 372
rect -557 332 -499 338
rect -365 372 -307 378
rect -365 338 -353 372
rect -319 338 -307 372
rect -365 332 -307 338
rect -173 372 -115 378
rect -173 338 -161 372
rect -127 338 -115 372
rect -173 332 -115 338
rect 19 372 77 378
rect 19 338 31 372
rect 65 338 77 372
rect 19 332 77 338
rect 211 372 269 378
rect 211 338 223 372
rect 257 338 269 372
rect 211 332 269 338
rect 403 372 461 378
rect 403 338 415 372
rect 449 338 461 372
rect 403 332 461 338
rect 595 372 653 378
rect 595 338 607 372
rect 641 338 653 372
rect 595 332 653 338
rect 787 372 845 378
rect 787 338 799 372
rect 833 338 845 372
rect 787 332 845 338
rect 979 372 1037 378
rect 979 338 991 372
rect 1025 338 1037 372
rect 979 332 1037 338
rect 1171 372 1229 378
rect 1171 338 1183 372
rect 1217 338 1229 372
rect 1171 332 1229 338
rect 1363 372 1421 378
rect 1363 338 1375 372
rect 1409 338 1421 372
rect 1363 332 1421 338
rect 1555 372 1613 378
rect 1555 338 1567 372
rect 1601 338 1613 372
rect 1555 332 1613 338
rect 1747 372 1805 378
rect 1747 338 1759 372
rect 1793 338 1805 372
rect 1747 332 1805 338
rect 1939 372 1997 378
rect 1939 338 1951 372
rect 1985 338 1997 372
rect 1939 332 1997 338
rect 2131 372 2189 378
rect 2131 338 2143 372
rect 2177 338 2189 372
rect 2131 332 2189 338
rect 2323 372 2381 378
rect 2323 338 2335 372
rect 2369 338 2381 372
rect 2323 332 2381 338
rect 2515 372 2573 378
rect 2515 338 2527 372
rect 2561 338 2573 372
rect 2515 332 2573 338
rect 2707 372 2765 378
rect 2707 338 2719 372
rect 2753 338 2765 372
rect 2707 332 2765 338
rect 2899 372 2957 378
rect 2899 338 2911 372
rect 2945 338 2957 372
rect 2899 332 2957 338
rect 3091 372 3149 378
rect 3091 338 3103 372
rect 3137 338 3149 372
rect 3091 332 3149 338
rect 3283 372 3341 378
rect 3283 338 3295 372
rect 3329 338 3341 372
rect 3283 332 3341 338
rect 3475 372 3533 378
rect 3475 338 3487 372
rect 3521 338 3533 372
rect 3475 332 3533 338
rect 3667 372 3725 378
rect 3667 338 3679 372
rect 3713 338 3725 372
rect 3667 332 3725 338
rect 3859 372 3917 378
rect 3859 338 3871 372
rect 3905 338 3917 372
rect 3859 332 3917 338
rect 4051 372 4109 378
rect 4051 338 4063 372
rect 4097 338 4109 372
rect 4051 332 4109 338
rect 4243 372 4301 378
rect 4243 338 4255 372
rect 4289 338 4301 372
rect 4243 332 4301 338
rect -4343 288 -4297 300
rect -4343 -288 -4337 288
rect -4303 -288 -4297 288
rect -4343 -300 -4297 -288
rect -4247 288 -4201 300
rect -4247 -288 -4241 288
rect -4207 -288 -4201 288
rect -4247 -300 -4201 -288
rect -4151 288 -4105 300
rect -4151 -288 -4145 288
rect -4111 -288 -4105 288
rect -4151 -300 -4105 -288
rect -4055 288 -4009 300
rect -4055 -288 -4049 288
rect -4015 -288 -4009 288
rect -4055 -300 -4009 -288
rect -3959 288 -3913 300
rect -3959 -288 -3953 288
rect -3919 -288 -3913 288
rect -3959 -300 -3913 -288
rect -3863 288 -3817 300
rect -3863 -288 -3857 288
rect -3823 -288 -3817 288
rect -3863 -300 -3817 -288
rect -3767 288 -3721 300
rect -3767 -288 -3761 288
rect -3727 -288 -3721 288
rect -3767 -300 -3721 -288
rect -3671 288 -3625 300
rect -3671 -288 -3665 288
rect -3631 -288 -3625 288
rect -3671 -300 -3625 -288
rect -3575 288 -3529 300
rect -3575 -288 -3569 288
rect -3535 -288 -3529 288
rect -3575 -300 -3529 -288
rect -3479 288 -3433 300
rect -3479 -288 -3473 288
rect -3439 -288 -3433 288
rect -3479 -300 -3433 -288
rect -3383 288 -3337 300
rect -3383 -288 -3377 288
rect -3343 -288 -3337 288
rect -3383 -300 -3337 -288
rect -3287 288 -3241 300
rect -3287 -288 -3281 288
rect -3247 -288 -3241 288
rect -3287 -300 -3241 -288
rect -3191 288 -3145 300
rect -3191 -288 -3185 288
rect -3151 -288 -3145 288
rect -3191 -300 -3145 -288
rect -3095 288 -3049 300
rect -3095 -288 -3089 288
rect -3055 -288 -3049 288
rect -3095 -300 -3049 -288
rect -2999 288 -2953 300
rect -2999 -288 -2993 288
rect -2959 -288 -2953 288
rect -2999 -300 -2953 -288
rect -2903 288 -2857 300
rect -2903 -288 -2897 288
rect -2863 -288 -2857 288
rect -2903 -300 -2857 -288
rect -2807 288 -2761 300
rect -2807 -288 -2801 288
rect -2767 -288 -2761 288
rect -2807 -300 -2761 -288
rect -2711 288 -2665 300
rect -2711 -288 -2705 288
rect -2671 -288 -2665 288
rect -2711 -300 -2665 -288
rect -2615 288 -2569 300
rect -2615 -288 -2609 288
rect -2575 -288 -2569 288
rect -2615 -300 -2569 -288
rect -2519 288 -2473 300
rect -2519 -288 -2513 288
rect -2479 -288 -2473 288
rect -2519 -300 -2473 -288
rect -2423 288 -2377 300
rect -2423 -288 -2417 288
rect -2383 -288 -2377 288
rect -2423 -300 -2377 -288
rect -2327 288 -2281 300
rect -2327 -288 -2321 288
rect -2287 -288 -2281 288
rect -2327 -300 -2281 -288
rect -2231 288 -2185 300
rect -2231 -288 -2225 288
rect -2191 -288 -2185 288
rect -2231 -300 -2185 -288
rect -2135 288 -2089 300
rect -2135 -288 -2129 288
rect -2095 -288 -2089 288
rect -2135 -300 -2089 -288
rect -2039 288 -1993 300
rect -2039 -288 -2033 288
rect -1999 -288 -1993 288
rect -2039 -300 -1993 -288
rect -1943 288 -1897 300
rect -1943 -288 -1937 288
rect -1903 -288 -1897 288
rect -1943 -300 -1897 -288
rect -1847 288 -1801 300
rect -1847 -288 -1841 288
rect -1807 -288 -1801 288
rect -1847 -300 -1801 -288
rect -1751 288 -1705 300
rect -1751 -288 -1745 288
rect -1711 -288 -1705 288
rect -1751 -300 -1705 -288
rect -1655 288 -1609 300
rect -1655 -288 -1649 288
rect -1615 -288 -1609 288
rect -1655 -300 -1609 -288
rect -1559 288 -1513 300
rect -1559 -288 -1553 288
rect -1519 -288 -1513 288
rect -1559 -300 -1513 -288
rect -1463 288 -1417 300
rect -1463 -288 -1457 288
rect -1423 -288 -1417 288
rect -1463 -300 -1417 -288
rect -1367 288 -1321 300
rect -1367 -288 -1361 288
rect -1327 -288 -1321 288
rect -1367 -300 -1321 -288
rect -1271 288 -1225 300
rect -1271 -288 -1265 288
rect -1231 -288 -1225 288
rect -1271 -300 -1225 -288
rect -1175 288 -1129 300
rect -1175 -288 -1169 288
rect -1135 -288 -1129 288
rect -1175 -300 -1129 -288
rect -1079 288 -1033 300
rect -1079 -288 -1073 288
rect -1039 -288 -1033 288
rect -1079 -300 -1033 -288
rect -983 288 -937 300
rect -983 -288 -977 288
rect -943 -288 -937 288
rect -983 -300 -937 -288
rect -887 288 -841 300
rect -887 -288 -881 288
rect -847 -288 -841 288
rect -887 -300 -841 -288
rect -791 288 -745 300
rect -791 -288 -785 288
rect -751 -288 -745 288
rect -791 -300 -745 -288
rect -695 288 -649 300
rect -695 -288 -689 288
rect -655 -288 -649 288
rect -695 -300 -649 -288
rect -599 288 -553 300
rect -599 -288 -593 288
rect -559 -288 -553 288
rect -599 -300 -553 -288
rect -503 288 -457 300
rect -503 -288 -497 288
rect -463 -288 -457 288
rect -503 -300 -457 -288
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect 457 288 503 300
rect 457 -288 463 288
rect 497 -288 503 288
rect 457 -300 503 -288
rect 553 288 599 300
rect 553 -288 559 288
rect 593 -288 599 288
rect 553 -300 599 -288
rect 649 288 695 300
rect 649 -288 655 288
rect 689 -288 695 288
rect 649 -300 695 -288
rect 745 288 791 300
rect 745 -288 751 288
rect 785 -288 791 288
rect 745 -300 791 -288
rect 841 288 887 300
rect 841 -288 847 288
rect 881 -288 887 288
rect 841 -300 887 -288
rect 937 288 983 300
rect 937 -288 943 288
rect 977 -288 983 288
rect 937 -300 983 -288
rect 1033 288 1079 300
rect 1033 -288 1039 288
rect 1073 -288 1079 288
rect 1033 -300 1079 -288
rect 1129 288 1175 300
rect 1129 -288 1135 288
rect 1169 -288 1175 288
rect 1129 -300 1175 -288
rect 1225 288 1271 300
rect 1225 -288 1231 288
rect 1265 -288 1271 288
rect 1225 -300 1271 -288
rect 1321 288 1367 300
rect 1321 -288 1327 288
rect 1361 -288 1367 288
rect 1321 -300 1367 -288
rect 1417 288 1463 300
rect 1417 -288 1423 288
rect 1457 -288 1463 288
rect 1417 -300 1463 -288
rect 1513 288 1559 300
rect 1513 -288 1519 288
rect 1553 -288 1559 288
rect 1513 -300 1559 -288
rect 1609 288 1655 300
rect 1609 -288 1615 288
rect 1649 -288 1655 288
rect 1609 -300 1655 -288
rect 1705 288 1751 300
rect 1705 -288 1711 288
rect 1745 -288 1751 288
rect 1705 -300 1751 -288
rect 1801 288 1847 300
rect 1801 -288 1807 288
rect 1841 -288 1847 288
rect 1801 -300 1847 -288
rect 1897 288 1943 300
rect 1897 -288 1903 288
rect 1937 -288 1943 288
rect 1897 -300 1943 -288
rect 1993 288 2039 300
rect 1993 -288 1999 288
rect 2033 -288 2039 288
rect 1993 -300 2039 -288
rect 2089 288 2135 300
rect 2089 -288 2095 288
rect 2129 -288 2135 288
rect 2089 -300 2135 -288
rect 2185 288 2231 300
rect 2185 -288 2191 288
rect 2225 -288 2231 288
rect 2185 -300 2231 -288
rect 2281 288 2327 300
rect 2281 -288 2287 288
rect 2321 -288 2327 288
rect 2281 -300 2327 -288
rect 2377 288 2423 300
rect 2377 -288 2383 288
rect 2417 -288 2423 288
rect 2377 -300 2423 -288
rect 2473 288 2519 300
rect 2473 -288 2479 288
rect 2513 -288 2519 288
rect 2473 -300 2519 -288
rect 2569 288 2615 300
rect 2569 -288 2575 288
rect 2609 -288 2615 288
rect 2569 -300 2615 -288
rect 2665 288 2711 300
rect 2665 -288 2671 288
rect 2705 -288 2711 288
rect 2665 -300 2711 -288
rect 2761 288 2807 300
rect 2761 -288 2767 288
rect 2801 -288 2807 288
rect 2761 -300 2807 -288
rect 2857 288 2903 300
rect 2857 -288 2863 288
rect 2897 -288 2903 288
rect 2857 -300 2903 -288
rect 2953 288 2999 300
rect 2953 -288 2959 288
rect 2993 -288 2999 288
rect 2953 -300 2999 -288
rect 3049 288 3095 300
rect 3049 -288 3055 288
rect 3089 -288 3095 288
rect 3049 -300 3095 -288
rect 3145 288 3191 300
rect 3145 -288 3151 288
rect 3185 -288 3191 288
rect 3145 -300 3191 -288
rect 3241 288 3287 300
rect 3241 -288 3247 288
rect 3281 -288 3287 288
rect 3241 -300 3287 -288
rect 3337 288 3383 300
rect 3337 -288 3343 288
rect 3377 -288 3383 288
rect 3337 -300 3383 -288
rect 3433 288 3479 300
rect 3433 -288 3439 288
rect 3473 -288 3479 288
rect 3433 -300 3479 -288
rect 3529 288 3575 300
rect 3529 -288 3535 288
rect 3569 -288 3575 288
rect 3529 -300 3575 -288
rect 3625 288 3671 300
rect 3625 -288 3631 288
rect 3665 -288 3671 288
rect 3625 -300 3671 -288
rect 3721 288 3767 300
rect 3721 -288 3727 288
rect 3761 -288 3767 288
rect 3721 -300 3767 -288
rect 3817 288 3863 300
rect 3817 -288 3823 288
rect 3857 -288 3863 288
rect 3817 -300 3863 -288
rect 3913 288 3959 300
rect 3913 -288 3919 288
rect 3953 -288 3959 288
rect 3913 -300 3959 -288
rect 4009 288 4055 300
rect 4009 -288 4015 288
rect 4049 -288 4055 288
rect 4009 -300 4055 -288
rect 4105 288 4151 300
rect 4105 -288 4111 288
rect 4145 -288 4151 288
rect 4105 -300 4151 -288
rect 4201 288 4247 300
rect 4201 -288 4207 288
rect 4241 -288 4247 288
rect 4201 -300 4247 -288
rect 4297 288 4343 300
rect 4297 -288 4303 288
rect 4337 -288 4343 288
rect 4297 -300 4343 -288
rect -4301 -338 -4243 -332
rect -4301 -372 -4289 -338
rect -4255 -372 -4243 -338
rect -4301 -378 -4243 -372
rect -4109 -338 -4051 -332
rect -4109 -372 -4097 -338
rect -4063 -372 -4051 -338
rect -4109 -378 -4051 -372
rect -3917 -338 -3859 -332
rect -3917 -372 -3905 -338
rect -3871 -372 -3859 -338
rect -3917 -378 -3859 -372
rect -3725 -338 -3667 -332
rect -3725 -372 -3713 -338
rect -3679 -372 -3667 -338
rect -3725 -378 -3667 -372
rect -3533 -338 -3475 -332
rect -3533 -372 -3521 -338
rect -3487 -372 -3475 -338
rect -3533 -378 -3475 -372
rect -3341 -338 -3283 -332
rect -3341 -372 -3329 -338
rect -3295 -372 -3283 -338
rect -3341 -378 -3283 -372
rect -3149 -338 -3091 -332
rect -3149 -372 -3137 -338
rect -3103 -372 -3091 -338
rect -3149 -378 -3091 -372
rect -2957 -338 -2899 -332
rect -2957 -372 -2945 -338
rect -2911 -372 -2899 -338
rect -2957 -378 -2899 -372
rect -2765 -338 -2707 -332
rect -2765 -372 -2753 -338
rect -2719 -372 -2707 -338
rect -2765 -378 -2707 -372
rect -2573 -338 -2515 -332
rect -2573 -372 -2561 -338
rect -2527 -372 -2515 -338
rect -2573 -378 -2515 -372
rect -2381 -338 -2323 -332
rect -2381 -372 -2369 -338
rect -2335 -372 -2323 -338
rect -2381 -378 -2323 -372
rect -2189 -338 -2131 -332
rect -2189 -372 -2177 -338
rect -2143 -372 -2131 -338
rect -2189 -378 -2131 -372
rect -1997 -338 -1939 -332
rect -1997 -372 -1985 -338
rect -1951 -372 -1939 -338
rect -1997 -378 -1939 -372
rect -1805 -338 -1747 -332
rect -1805 -372 -1793 -338
rect -1759 -372 -1747 -338
rect -1805 -378 -1747 -372
rect -1613 -338 -1555 -332
rect -1613 -372 -1601 -338
rect -1567 -372 -1555 -338
rect -1613 -378 -1555 -372
rect -1421 -338 -1363 -332
rect -1421 -372 -1409 -338
rect -1375 -372 -1363 -338
rect -1421 -378 -1363 -372
rect -1229 -338 -1171 -332
rect -1229 -372 -1217 -338
rect -1183 -372 -1171 -338
rect -1229 -378 -1171 -372
rect -1037 -338 -979 -332
rect -1037 -372 -1025 -338
rect -991 -372 -979 -338
rect -1037 -378 -979 -372
rect -845 -338 -787 -332
rect -845 -372 -833 -338
rect -799 -372 -787 -338
rect -845 -378 -787 -372
rect -653 -338 -595 -332
rect -653 -372 -641 -338
rect -607 -372 -595 -338
rect -653 -378 -595 -372
rect -461 -338 -403 -332
rect -461 -372 -449 -338
rect -415 -372 -403 -338
rect -461 -378 -403 -372
rect -269 -338 -211 -332
rect -269 -372 -257 -338
rect -223 -372 -211 -338
rect -269 -378 -211 -372
rect -77 -338 -19 -332
rect -77 -372 -65 -338
rect -31 -372 -19 -338
rect -77 -378 -19 -372
rect 115 -338 173 -332
rect 115 -372 127 -338
rect 161 -372 173 -338
rect 115 -378 173 -372
rect 307 -338 365 -332
rect 307 -372 319 -338
rect 353 -372 365 -338
rect 307 -378 365 -372
rect 499 -338 557 -332
rect 499 -372 511 -338
rect 545 -372 557 -338
rect 499 -378 557 -372
rect 691 -338 749 -332
rect 691 -372 703 -338
rect 737 -372 749 -338
rect 691 -378 749 -372
rect 883 -338 941 -332
rect 883 -372 895 -338
rect 929 -372 941 -338
rect 883 -378 941 -372
rect 1075 -338 1133 -332
rect 1075 -372 1087 -338
rect 1121 -372 1133 -338
rect 1075 -378 1133 -372
rect 1267 -338 1325 -332
rect 1267 -372 1279 -338
rect 1313 -372 1325 -338
rect 1267 -378 1325 -372
rect 1459 -338 1517 -332
rect 1459 -372 1471 -338
rect 1505 -372 1517 -338
rect 1459 -378 1517 -372
rect 1651 -338 1709 -332
rect 1651 -372 1663 -338
rect 1697 -372 1709 -338
rect 1651 -378 1709 -372
rect 1843 -338 1901 -332
rect 1843 -372 1855 -338
rect 1889 -372 1901 -338
rect 1843 -378 1901 -372
rect 2035 -338 2093 -332
rect 2035 -372 2047 -338
rect 2081 -372 2093 -338
rect 2035 -378 2093 -372
rect 2227 -338 2285 -332
rect 2227 -372 2239 -338
rect 2273 -372 2285 -338
rect 2227 -378 2285 -372
rect 2419 -338 2477 -332
rect 2419 -372 2431 -338
rect 2465 -372 2477 -338
rect 2419 -378 2477 -372
rect 2611 -338 2669 -332
rect 2611 -372 2623 -338
rect 2657 -372 2669 -338
rect 2611 -378 2669 -372
rect 2803 -338 2861 -332
rect 2803 -372 2815 -338
rect 2849 -372 2861 -338
rect 2803 -378 2861 -372
rect 2995 -338 3053 -332
rect 2995 -372 3007 -338
rect 3041 -372 3053 -338
rect 2995 -378 3053 -372
rect 3187 -338 3245 -332
rect 3187 -372 3199 -338
rect 3233 -372 3245 -338
rect 3187 -378 3245 -372
rect 3379 -338 3437 -332
rect 3379 -372 3391 -338
rect 3425 -372 3437 -338
rect 3379 -378 3437 -372
rect 3571 -338 3629 -332
rect 3571 -372 3583 -338
rect 3617 -372 3629 -338
rect 3571 -378 3629 -372
rect 3763 -338 3821 -332
rect 3763 -372 3775 -338
rect 3809 -372 3821 -338
rect 3763 -378 3821 -372
rect 3955 -338 4013 -332
rect 3955 -372 3967 -338
rect 4001 -372 4013 -338
rect 3955 -378 4013 -372
rect 4147 -338 4205 -332
rect 4147 -372 4159 -338
rect 4193 -372 4205 -338
rect 4147 -378 4205 -372
<< properties >>
string FIXED_BBOX -4434 -457 4434 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 90 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
