magic
tech sky130A
magscale 1 2
timestamp 1707380652
<< error_s >>
rect 438 870 468 879
rect 434 824 476 835
rect 400 790 510 801
rect 1987 670 2021 678
rect 176 614 218 648
rect 2006 634 2040 644
rect 2006 620 2016 634
rect 2030 620 2040 634
rect 176 604 222 614
rect 2006 610 2040 620
rect 210 570 244 580
<< polycont >>
rect 2006 610 2040 644
rect 1904 -104 1938 -70
rect 1978 -646 2012 -612
<< locali >>
rect 218 604 222 648
rect 1356 -64 1780 -58
rect 1356 -104 1712 -64
rect 1432 -106 1712 -104
rect 1774 -106 1780 -64
<< viali >>
rect 434 824 476 870
rect 176 604 218 648
rect 2002 644 2046 646
rect 2002 610 2006 644
rect 2006 610 2040 644
rect 2040 610 2046 644
rect 2002 606 2046 610
rect 2256 -34 2316 16
rect 984 -104 1032 -60
rect 1712 -106 1774 -64
rect 1892 -70 1936 -66
rect 1892 -102 1904 -70
rect 1904 -102 1936 -70
rect 2070 -100 2128 -58
rect 142 -652 188 -610
rect 1962 -612 2012 -606
rect 1962 -646 1978 -612
rect 1978 -646 2012 -612
rect 1962 -652 2012 -646
rect 410 -884 456 -848
<< metal1 >>
rect -292 978 -92 982
rect -292 906 -230 978
rect -158 906 -92 978
rect 152 910 162 982
rect 234 910 244 982
rect -292 782 -92 906
rect 420 870 488 916
rect 2112 894 2674 984
rect 420 824 434 870
rect 476 824 488 870
rect 420 820 488 824
rect 428 812 482 820
rect -580 652 -338 690
rect -580 568 -504 652
rect -402 568 -338 652
rect 158 594 168 658
rect 226 594 236 658
rect 1990 646 2058 652
rect 1990 606 2002 646
rect 2046 644 2058 646
rect 2046 606 2460 644
rect 1990 600 2058 606
rect -580 462 -338 568
rect 722 528 732 592
rect 804 542 914 592
rect 2402 572 2452 606
rect 804 528 846 542
rect 2384 516 2394 572
rect 2456 516 2466 572
rect -276 -358 -76 -250
rect -276 -430 -232 -358
rect -152 -430 -76 -358
rect -276 -450 -76 -430
rect 120 -432 130 -360
rect 210 -432 220 -360
rect 334 -436 414 444
rect 1326 200 1852 256
rect 2238 190 2248 262
rect 2326 190 2336 262
rect 2244 16 2328 22
rect 2402 16 2452 516
rect 2570 266 2660 894
rect 2756 572 2956 650
rect 2756 512 2830 572
rect 2898 512 2956 572
rect 2756 450 2956 512
rect 2564 194 2574 266
rect 2652 194 2662 266
rect 2242 -34 2256 16
rect 2316 -34 2452 16
rect 2242 -36 2452 -34
rect 2244 -40 2328 -36
rect 972 -60 1044 -54
rect 2058 -58 2140 -52
rect 956 -112 966 -60
rect 1040 -112 1050 -60
rect 1700 -62 1786 -58
rect 1880 -62 1948 -60
rect 1700 -64 1948 -62
rect 1700 -106 1712 -64
rect 1774 -66 1948 -64
rect 1774 -102 1892 -66
rect 1936 -102 1948 -66
rect 1774 -104 1948 -102
rect 1774 -106 1786 -104
rect 1700 -112 1786 -106
rect 1880 -108 1948 -104
rect 2058 -100 2070 -58
rect 2128 -100 2140 -58
rect 2058 -106 2140 -100
rect 2078 -136 2128 -106
rect 2078 -140 2442 -136
rect 2078 -180 2444 -140
rect 2388 -464 2444 -180
rect 2372 -524 2382 -464
rect 2450 -524 2460 -464
rect -600 -590 -400 -538
rect -600 -688 -568 -590
rect -456 -688 -400 -590
rect 874 -592 884 -534
rect 940 -592 950 -534
rect 2388 -596 2444 -524
rect 2370 -598 2444 -596
rect 1956 -600 2444 -598
rect 110 -660 120 -602
rect 194 -660 204 -602
rect 1950 -606 2444 -600
rect 1950 -652 1962 -606
rect 2012 -642 2444 -606
rect 2012 -652 2430 -642
rect 1950 -654 2430 -652
rect 1950 -656 2370 -654
rect 1950 -658 2024 -656
rect -600 -738 -400 -688
rect 398 -848 468 -842
rect 398 -884 410 -848
rect 456 -884 468 -848
rect 398 -916 468 -884
rect 2570 -894 2660 194
rect 2766 -452 2966 -368
rect 2766 -512 2822 -452
rect 2890 -512 2966 -452
rect 2766 -568 2966 -512
rect 2076 -980 2660 -894
rect 2076 -984 2638 -980
<< via1 >>
rect -230 906 -158 978
rect 162 910 234 982
rect -504 568 -402 652
rect 168 648 226 658
rect 168 604 176 648
rect 176 604 218 648
rect 218 604 226 648
rect 168 594 226 604
rect 732 528 804 592
rect 2394 516 2456 572
rect -232 -430 -152 -358
rect 130 -432 210 -360
rect 2248 190 2326 262
rect 2830 512 2898 572
rect 2574 194 2652 266
rect 966 -104 984 -60
rect 984 -104 1032 -60
rect 1032 -104 1040 -60
rect 966 -112 1040 -104
rect 2382 -524 2450 -464
rect -568 -688 -456 -590
rect 884 -592 940 -534
rect 120 -610 194 -602
rect 120 -652 142 -610
rect 142 -652 188 -610
rect 188 -652 194 -610
rect 120 -660 194 -652
rect 2822 -512 2890 -452
<< metal2 >>
rect -230 984 -158 988
rect 162 984 234 992
rect -234 982 238 984
rect -234 978 162 982
rect -234 908 -230 978
rect -158 910 162 978
rect 234 910 238 982
rect -158 908 238 910
rect -230 896 -158 906
rect 162 900 234 908
rect -504 656 -402 662
rect 168 658 226 668
rect -504 652 168 656
rect -402 610 168 652
rect 168 584 226 594
rect 732 592 804 602
rect -504 558 -402 568
rect 2394 572 2456 582
rect 2830 572 2898 582
rect 804 528 808 542
rect 732 486 808 528
rect 2392 516 2394 572
rect 2456 516 2830 572
rect 2392 514 2830 516
rect 2394 506 2456 514
rect 2898 514 2902 572
rect 2830 502 2898 512
rect 732 -56 798 486
rect 2248 266 2326 272
rect 2574 266 2652 276
rect 2244 262 2574 266
rect 2244 194 2248 262
rect 2326 194 2574 262
rect 2248 180 2326 190
rect 2574 184 2652 194
rect 966 -56 1040 -50
rect 730 -60 1040 -56
rect 730 -112 966 -60
rect 730 -116 1040 -112
rect -232 -358 -152 -348
rect 130 -360 210 -350
rect -152 -430 130 -364
rect -232 -432 130 -430
rect -232 -434 210 -432
rect -232 -440 -152 -434
rect 130 -442 210 -434
rect 732 -494 798 -116
rect 966 -122 1040 -116
rect 2822 -452 2890 -442
rect 2382 -464 2450 -454
rect 732 -534 940 -494
rect 2372 -518 2382 -464
rect 2450 -512 2822 -464
rect 2450 -518 2890 -512
rect 2822 -522 2890 -518
rect 2382 -534 2450 -524
rect -568 -590 -456 -580
rect 734 -592 884 -534
rect 940 -592 962 -534
rect 120 -596 194 -592
rect -456 -602 194 -596
rect 884 -594 962 -592
rect 884 -602 940 -594
rect -456 -660 120 -602
rect -456 -664 194 -660
rect 120 -670 194 -664
rect -568 -698 -456 -688
use sky130_fd_sc_hd__dfrbp_2  sky130_fd_sc_hd__dfrbp_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 2362 0 1 394
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 2334 0 1 -320
box -38 -48 590 592
use sky130_fd_sc_hd__dfrbp_2  x3
timestamp 1705271942
transform 1 0 124 0 -1 -396
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform -1 0 1418 0 1 -320
box -38 -48 498 592
<< labels >>
flabel metal1 2766 -568 2966 -368 0 FreeSans 256 0 0 0 QB
port 4 nsew
flabel metal1 2756 450 2956 650 0 FreeSans 256 0 0 0 QA
port 3 nsew
flabel metal1 -600 -738 -400 -538 0 FreeSans 256 0 0 0 B
port 5 nsew
flabel metal1 -276 -450 -76 -250 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 -580 462 -338 690 0 FreeSans 256 0 0 0 A
port 6 nsew
flabel metal1 -292 782 -92 982 0 FreeSans 256 0 0 0 VDD
port 1 nsew
<< end >>
