** sch_path: /home/harsh/design/xschem/inverter.sch
.subckt inverter inp out VDD VSS
*.PININFO inp:I out:O VDD:B VSS:B
x4 inp VSS VSS VDD VDD out sky130_fd_sc_hd__inv_4
.ends
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.end
