magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -1325 881 -1267 887
rect -1133 881 -1075 887
rect -941 881 -883 887
rect -749 881 -691 887
rect -557 881 -499 887
rect -365 881 -307 887
rect -173 881 -115 887
rect 19 881 77 887
rect 211 881 269 887
rect 403 881 461 887
rect 595 881 653 887
rect 787 881 845 887
rect 979 881 1037 887
rect 1171 881 1229 887
rect 1363 881 1421 887
rect -1325 847 -1313 881
rect -1133 847 -1121 881
rect -941 847 -929 881
rect -749 847 -737 881
rect -557 847 -545 881
rect -365 847 -353 881
rect -173 847 -161 881
rect 19 847 31 881
rect 211 847 223 881
rect 403 847 415 881
rect 595 847 607 881
rect 787 847 799 881
rect 979 847 991 881
rect 1171 847 1183 881
rect 1363 847 1375 881
rect -1325 841 -1267 847
rect -1133 841 -1075 847
rect -941 841 -883 847
rect -749 841 -691 847
rect -557 841 -499 847
rect -365 841 -307 847
rect -173 841 -115 847
rect 19 841 77 847
rect 211 841 269 847
rect 403 841 461 847
rect 595 841 653 847
rect 787 841 845 847
rect 979 841 1037 847
rect 1171 841 1229 847
rect 1363 841 1421 847
rect -1421 -847 -1363 -841
rect -1229 -847 -1171 -841
rect -1037 -847 -979 -841
rect -845 -847 -787 -841
rect -653 -847 -595 -841
rect -461 -847 -403 -841
rect -269 -847 -211 -841
rect -77 -847 -19 -841
rect 115 -847 173 -841
rect 307 -847 365 -841
rect 499 -847 557 -841
rect 691 -847 749 -841
rect 883 -847 941 -841
rect 1075 -847 1133 -841
rect 1267 -847 1325 -841
rect -1421 -881 -1409 -847
rect -1229 -881 -1217 -847
rect -1037 -881 -1025 -847
rect -845 -881 -833 -847
rect -653 -881 -641 -847
rect -461 -881 -449 -847
rect -269 -881 -257 -847
rect -77 -881 -65 -847
rect 115 -881 127 -847
rect 307 -881 319 -847
rect 499 -881 511 -847
rect 691 -881 703 -847
rect 883 -881 895 -847
rect 1075 -881 1087 -847
rect 1267 -881 1279 -847
rect -1421 -887 -1363 -881
rect -1229 -887 -1171 -881
rect -1037 -887 -979 -881
rect -845 -887 -787 -881
rect -653 -887 -595 -881
rect -461 -887 -403 -881
rect -269 -887 -211 -881
rect -77 -887 -19 -881
rect 115 -887 173 -881
rect 307 -887 365 -881
rect 499 -887 557 -881
rect 691 -887 749 -881
rect 883 -887 941 -881
rect 1075 -887 1133 -881
rect 1267 -887 1325 -881
<< nwell >>
rect -1607 -1019 1607 1019
<< pmos >>
rect -1407 -800 -1377 800
rect -1311 -800 -1281 800
rect -1215 -800 -1185 800
rect -1119 -800 -1089 800
rect -1023 -800 -993 800
rect -927 -800 -897 800
rect -831 -800 -801 800
rect -735 -800 -705 800
rect -639 -800 -609 800
rect -543 -800 -513 800
rect -447 -800 -417 800
rect -351 -800 -321 800
rect -255 -800 -225 800
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
rect 225 -800 255 800
rect 321 -800 351 800
rect 417 -800 447 800
rect 513 -800 543 800
rect 609 -800 639 800
rect 705 -800 735 800
rect 801 -800 831 800
rect 897 -800 927 800
rect 993 -800 1023 800
rect 1089 -800 1119 800
rect 1185 -800 1215 800
rect 1281 -800 1311 800
rect 1377 -800 1407 800
<< pdiff >>
rect -1469 788 -1407 800
rect -1469 -788 -1457 788
rect -1423 -788 -1407 788
rect -1469 -800 -1407 -788
rect -1377 788 -1311 800
rect -1377 -788 -1361 788
rect -1327 -788 -1311 788
rect -1377 -800 -1311 -788
rect -1281 788 -1215 800
rect -1281 -788 -1265 788
rect -1231 -788 -1215 788
rect -1281 -800 -1215 -788
rect -1185 788 -1119 800
rect -1185 -788 -1169 788
rect -1135 -788 -1119 788
rect -1185 -800 -1119 -788
rect -1089 788 -1023 800
rect -1089 -788 -1073 788
rect -1039 -788 -1023 788
rect -1089 -800 -1023 -788
rect -993 788 -927 800
rect -993 -788 -977 788
rect -943 -788 -927 788
rect -993 -800 -927 -788
rect -897 788 -831 800
rect -897 -788 -881 788
rect -847 -788 -831 788
rect -897 -800 -831 -788
rect -801 788 -735 800
rect -801 -788 -785 788
rect -751 -788 -735 788
rect -801 -800 -735 -788
rect -705 788 -639 800
rect -705 -788 -689 788
rect -655 -788 -639 788
rect -705 -800 -639 -788
rect -609 788 -543 800
rect -609 -788 -593 788
rect -559 -788 -543 788
rect -609 -800 -543 -788
rect -513 788 -447 800
rect -513 -788 -497 788
rect -463 -788 -447 788
rect -513 -800 -447 -788
rect -417 788 -351 800
rect -417 -788 -401 788
rect -367 -788 -351 788
rect -417 -800 -351 -788
rect -321 788 -255 800
rect -321 -788 -305 788
rect -271 -788 -255 788
rect -321 -800 -255 -788
rect -225 788 -159 800
rect -225 -788 -209 788
rect -175 -788 -159 788
rect -225 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 225 800
rect 159 -788 175 788
rect 209 -788 225 788
rect 159 -800 225 -788
rect 255 788 321 800
rect 255 -788 271 788
rect 305 -788 321 788
rect 255 -800 321 -788
rect 351 788 417 800
rect 351 -788 367 788
rect 401 -788 417 788
rect 351 -800 417 -788
rect 447 788 513 800
rect 447 -788 463 788
rect 497 -788 513 788
rect 447 -800 513 -788
rect 543 788 609 800
rect 543 -788 559 788
rect 593 -788 609 788
rect 543 -800 609 -788
rect 639 788 705 800
rect 639 -788 655 788
rect 689 -788 705 788
rect 639 -800 705 -788
rect 735 788 801 800
rect 735 -788 751 788
rect 785 -788 801 788
rect 735 -800 801 -788
rect 831 788 897 800
rect 831 -788 847 788
rect 881 -788 897 788
rect 831 -800 897 -788
rect 927 788 993 800
rect 927 -788 943 788
rect 977 -788 993 788
rect 927 -800 993 -788
rect 1023 788 1089 800
rect 1023 -788 1039 788
rect 1073 -788 1089 788
rect 1023 -800 1089 -788
rect 1119 788 1185 800
rect 1119 -788 1135 788
rect 1169 -788 1185 788
rect 1119 -800 1185 -788
rect 1215 788 1281 800
rect 1215 -788 1231 788
rect 1265 -788 1281 788
rect 1215 -800 1281 -788
rect 1311 788 1377 800
rect 1311 -788 1327 788
rect 1361 -788 1377 788
rect 1311 -800 1377 -788
rect 1407 788 1469 800
rect 1407 -788 1423 788
rect 1457 -788 1469 788
rect 1407 -800 1469 -788
<< pdiffc >>
rect -1457 -788 -1423 788
rect -1361 -788 -1327 788
rect -1265 -788 -1231 788
rect -1169 -788 -1135 788
rect -1073 -788 -1039 788
rect -977 -788 -943 788
rect -881 -788 -847 788
rect -785 -788 -751 788
rect -689 -788 -655 788
rect -593 -788 -559 788
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect 559 -788 593 788
rect 655 -788 689 788
rect 751 -788 785 788
rect 847 -788 881 788
rect 943 -788 977 788
rect 1039 -788 1073 788
rect 1135 -788 1169 788
rect 1231 -788 1265 788
rect 1327 -788 1361 788
rect 1423 -788 1457 788
<< nsubdiff >>
rect -1571 949 -1475 983
rect 1475 949 1571 983
rect -1571 887 -1537 949
rect 1537 887 1571 949
rect -1571 -949 -1537 -887
rect 1537 -949 1571 -887
rect -1571 -983 -1475 -949
rect 1475 -983 1571 -949
<< nsubdiffcont >>
rect -1475 949 1475 983
rect -1571 -887 -1537 887
rect 1537 -887 1571 887
rect -1475 -983 1475 -949
<< poly >>
rect -1329 881 -1263 897
rect -1329 847 -1313 881
rect -1279 847 -1263 881
rect -1329 831 -1263 847
rect -1137 881 -1071 897
rect -1137 847 -1121 881
rect -1087 847 -1071 881
rect -1137 831 -1071 847
rect -945 881 -879 897
rect -945 847 -929 881
rect -895 847 -879 881
rect -945 831 -879 847
rect -753 881 -687 897
rect -753 847 -737 881
rect -703 847 -687 881
rect -753 831 -687 847
rect -561 881 -495 897
rect -561 847 -545 881
rect -511 847 -495 881
rect -561 831 -495 847
rect -369 881 -303 897
rect -369 847 -353 881
rect -319 847 -303 881
rect -369 831 -303 847
rect -177 881 -111 897
rect -177 847 -161 881
rect -127 847 -111 881
rect -177 831 -111 847
rect 15 881 81 897
rect 15 847 31 881
rect 65 847 81 881
rect 15 831 81 847
rect 207 881 273 897
rect 207 847 223 881
rect 257 847 273 881
rect 207 831 273 847
rect 399 881 465 897
rect 399 847 415 881
rect 449 847 465 881
rect 399 831 465 847
rect 591 881 657 897
rect 591 847 607 881
rect 641 847 657 881
rect 591 831 657 847
rect 783 881 849 897
rect 783 847 799 881
rect 833 847 849 881
rect 783 831 849 847
rect 975 881 1041 897
rect 975 847 991 881
rect 1025 847 1041 881
rect 975 831 1041 847
rect 1167 881 1233 897
rect 1167 847 1183 881
rect 1217 847 1233 881
rect 1167 831 1233 847
rect 1359 881 1425 897
rect 1359 847 1375 881
rect 1409 847 1425 881
rect 1359 831 1425 847
rect -1407 800 -1377 826
rect -1311 800 -1281 831
rect -1215 800 -1185 826
rect -1119 800 -1089 831
rect -1023 800 -993 826
rect -927 800 -897 831
rect -831 800 -801 826
rect -735 800 -705 831
rect -639 800 -609 826
rect -543 800 -513 831
rect -447 800 -417 826
rect -351 800 -321 831
rect -255 800 -225 826
rect -159 800 -129 831
rect -63 800 -33 826
rect 33 800 63 831
rect 129 800 159 826
rect 225 800 255 831
rect 321 800 351 826
rect 417 800 447 831
rect 513 800 543 826
rect 609 800 639 831
rect 705 800 735 826
rect 801 800 831 831
rect 897 800 927 826
rect 993 800 1023 831
rect 1089 800 1119 826
rect 1185 800 1215 831
rect 1281 800 1311 826
rect 1377 800 1407 831
rect -1407 -831 -1377 -800
rect -1311 -826 -1281 -800
rect -1215 -831 -1185 -800
rect -1119 -826 -1089 -800
rect -1023 -831 -993 -800
rect -927 -826 -897 -800
rect -831 -831 -801 -800
rect -735 -826 -705 -800
rect -639 -831 -609 -800
rect -543 -826 -513 -800
rect -447 -831 -417 -800
rect -351 -826 -321 -800
rect -255 -831 -225 -800
rect -159 -826 -129 -800
rect -63 -831 -33 -800
rect 33 -826 63 -800
rect 129 -831 159 -800
rect 225 -826 255 -800
rect 321 -831 351 -800
rect 417 -826 447 -800
rect 513 -831 543 -800
rect 609 -826 639 -800
rect 705 -831 735 -800
rect 801 -826 831 -800
rect 897 -831 927 -800
rect 993 -826 1023 -800
rect 1089 -831 1119 -800
rect 1185 -826 1215 -800
rect 1281 -831 1311 -800
rect 1377 -826 1407 -800
rect -1425 -847 -1359 -831
rect -1425 -881 -1409 -847
rect -1375 -881 -1359 -847
rect -1425 -897 -1359 -881
rect -1233 -847 -1167 -831
rect -1233 -881 -1217 -847
rect -1183 -881 -1167 -847
rect -1233 -897 -1167 -881
rect -1041 -847 -975 -831
rect -1041 -881 -1025 -847
rect -991 -881 -975 -847
rect -1041 -897 -975 -881
rect -849 -847 -783 -831
rect -849 -881 -833 -847
rect -799 -881 -783 -847
rect -849 -897 -783 -881
rect -657 -847 -591 -831
rect -657 -881 -641 -847
rect -607 -881 -591 -847
rect -657 -897 -591 -881
rect -465 -847 -399 -831
rect -465 -881 -449 -847
rect -415 -881 -399 -847
rect -465 -897 -399 -881
rect -273 -847 -207 -831
rect -273 -881 -257 -847
rect -223 -881 -207 -847
rect -273 -897 -207 -881
rect -81 -847 -15 -831
rect -81 -881 -65 -847
rect -31 -881 -15 -847
rect -81 -897 -15 -881
rect 111 -847 177 -831
rect 111 -881 127 -847
rect 161 -881 177 -847
rect 111 -897 177 -881
rect 303 -847 369 -831
rect 303 -881 319 -847
rect 353 -881 369 -847
rect 303 -897 369 -881
rect 495 -847 561 -831
rect 495 -881 511 -847
rect 545 -881 561 -847
rect 495 -897 561 -881
rect 687 -847 753 -831
rect 687 -881 703 -847
rect 737 -881 753 -847
rect 687 -897 753 -881
rect 879 -847 945 -831
rect 879 -881 895 -847
rect 929 -881 945 -847
rect 879 -897 945 -881
rect 1071 -847 1137 -831
rect 1071 -881 1087 -847
rect 1121 -881 1137 -847
rect 1071 -897 1137 -881
rect 1263 -847 1329 -831
rect 1263 -881 1279 -847
rect 1313 -881 1329 -847
rect 1263 -897 1329 -881
<< polycont >>
rect -1313 847 -1279 881
rect -1121 847 -1087 881
rect -929 847 -895 881
rect -737 847 -703 881
rect -545 847 -511 881
rect -353 847 -319 881
rect -161 847 -127 881
rect 31 847 65 881
rect 223 847 257 881
rect 415 847 449 881
rect 607 847 641 881
rect 799 847 833 881
rect 991 847 1025 881
rect 1183 847 1217 881
rect 1375 847 1409 881
rect -1409 -881 -1375 -847
rect -1217 -881 -1183 -847
rect -1025 -881 -991 -847
rect -833 -881 -799 -847
rect -641 -881 -607 -847
rect -449 -881 -415 -847
rect -257 -881 -223 -847
rect -65 -881 -31 -847
rect 127 -881 161 -847
rect 319 -881 353 -847
rect 511 -881 545 -847
rect 703 -881 737 -847
rect 895 -881 929 -847
rect 1087 -881 1121 -847
rect 1279 -881 1313 -847
<< locali >>
rect -1571 949 -1475 983
rect 1475 949 1571 983
rect -1571 887 -1537 949
rect 1537 887 1571 949
rect -1329 847 -1313 881
rect -1279 847 -1263 881
rect -1137 847 -1121 881
rect -1087 847 -1071 881
rect -945 847 -929 881
rect -895 847 -879 881
rect -753 847 -737 881
rect -703 847 -687 881
rect -561 847 -545 881
rect -511 847 -495 881
rect -369 847 -353 881
rect -319 847 -303 881
rect -177 847 -161 881
rect -127 847 -111 881
rect 15 847 31 881
rect 65 847 81 881
rect 207 847 223 881
rect 257 847 273 881
rect 399 847 415 881
rect 449 847 465 881
rect 591 847 607 881
rect 641 847 657 881
rect 783 847 799 881
rect 833 847 849 881
rect 975 847 991 881
rect 1025 847 1041 881
rect 1167 847 1183 881
rect 1217 847 1233 881
rect 1359 847 1375 881
rect 1409 847 1425 881
rect -1457 788 -1423 804
rect -1457 -804 -1423 -788
rect -1361 788 -1327 804
rect -1361 -804 -1327 -788
rect -1265 788 -1231 804
rect -1265 -804 -1231 -788
rect -1169 788 -1135 804
rect -1169 -804 -1135 -788
rect -1073 788 -1039 804
rect -1073 -804 -1039 -788
rect -977 788 -943 804
rect -977 -804 -943 -788
rect -881 788 -847 804
rect -881 -804 -847 -788
rect -785 788 -751 804
rect -785 -804 -751 -788
rect -689 788 -655 804
rect -689 -804 -655 -788
rect -593 788 -559 804
rect -593 -804 -559 -788
rect -497 788 -463 804
rect -497 -804 -463 -788
rect -401 788 -367 804
rect -401 -804 -367 -788
rect -305 788 -271 804
rect -305 -804 -271 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 271 788 305 804
rect 271 -804 305 -788
rect 367 788 401 804
rect 367 -804 401 -788
rect 463 788 497 804
rect 463 -804 497 -788
rect 559 788 593 804
rect 559 -804 593 -788
rect 655 788 689 804
rect 655 -804 689 -788
rect 751 788 785 804
rect 751 -804 785 -788
rect 847 788 881 804
rect 847 -804 881 -788
rect 943 788 977 804
rect 943 -804 977 -788
rect 1039 788 1073 804
rect 1039 -804 1073 -788
rect 1135 788 1169 804
rect 1135 -804 1169 -788
rect 1231 788 1265 804
rect 1231 -804 1265 -788
rect 1327 788 1361 804
rect 1327 -804 1361 -788
rect 1423 788 1457 804
rect 1423 -804 1457 -788
rect -1425 -881 -1409 -847
rect -1375 -881 -1359 -847
rect -1233 -881 -1217 -847
rect -1183 -881 -1167 -847
rect -1041 -881 -1025 -847
rect -991 -881 -975 -847
rect -849 -881 -833 -847
rect -799 -881 -783 -847
rect -657 -881 -641 -847
rect -607 -881 -591 -847
rect -465 -881 -449 -847
rect -415 -881 -399 -847
rect -273 -881 -257 -847
rect -223 -881 -207 -847
rect -81 -881 -65 -847
rect -31 -881 -15 -847
rect 111 -881 127 -847
rect 161 -881 177 -847
rect 303 -881 319 -847
rect 353 -881 369 -847
rect 495 -881 511 -847
rect 545 -881 561 -847
rect 687 -881 703 -847
rect 737 -881 753 -847
rect 879 -881 895 -847
rect 929 -881 945 -847
rect 1071 -881 1087 -847
rect 1121 -881 1137 -847
rect 1263 -881 1279 -847
rect 1313 -881 1329 -847
rect -1571 -949 -1537 -887
rect 1537 -949 1571 -887
rect -1571 -983 -1475 -949
rect 1475 -983 1571 -949
<< viali >>
rect -1313 847 -1279 881
rect -1121 847 -1087 881
rect -929 847 -895 881
rect -737 847 -703 881
rect -545 847 -511 881
rect -353 847 -319 881
rect -161 847 -127 881
rect 31 847 65 881
rect 223 847 257 881
rect 415 847 449 881
rect 607 847 641 881
rect 799 847 833 881
rect 991 847 1025 881
rect 1183 847 1217 881
rect 1375 847 1409 881
rect -1457 -788 -1423 788
rect -1361 -788 -1327 788
rect -1265 -788 -1231 788
rect -1169 -788 -1135 788
rect -1073 -788 -1039 788
rect -977 -788 -943 788
rect -881 -788 -847 788
rect -785 -788 -751 788
rect -689 -788 -655 788
rect -593 -788 -559 788
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect 559 -788 593 788
rect 655 -788 689 788
rect 751 -788 785 788
rect 847 -788 881 788
rect 943 -788 977 788
rect 1039 -788 1073 788
rect 1135 -788 1169 788
rect 1231 -788 1265 788
rect 1327 -788 1361 788
rect 1423 -788 1457 788
rect -1409 -881 -1375 -847
rect -1217 -881 -1183 -847
rect -1025 -881 -991 -847
rect -833 -881 -799 -847
rect -641 -881 -607 -847
rect -449 -881 -415 -847
rect -257 -881 -223 -847
rect -65 -881 -31 -847
rect 127 -881 161 -847
rect 319 -881 353 -847
rect 511 -881 545 -847
rect 703 -881 737 -847
rect 895 -881 929 -847
rect 1087 -881 1121 -847
rect 1279 -881 1313 -847
<< metal1 >>
rect -1325 881 -1267 887
rect -1325 847 -1313 881
rect -1279 847 -1267 881
rect -1325 841 -1267 847
rect -1133 881 -1075 887
rect -1133 847 -1121 881
rect -1087 847 -1075 881
rect -1133 841 -1075 847
rect -941 881 -883 887
rect -941 847 -929 881
rect -895 847 -883 881
rect -941 841 -883 847
rect -749 881 -691 887
rect -749 847 -737 881
rect -703 847 -691 881
rect -749 841 -691 847
rect -557 881 -499 887
rect -557 847 -545 881
rect -511 847 -499 881
rect -557 841 -499 847
rect -365 881 -307 887
rect -365 847 -353 881
rect -319 847 -307 881
rect -365 841 -307 847
rect -173 881 -115 887
rect -173 847 -161 881
rect -127 847 -115 881
rect -173 841 -115 847
rect 19 881 77 887
rect 19 847 31 881
rect 65 847 77 881
rect 19 841 77 847
rect 211 881 269 887
rect 211 847 223 881
rect 257 847 269 881
rect 211 841 269 847
rect 403 881 461 887
rect 403 847 415 881
rect 449 847 461 881
rect 403 841 461 847
rect 595 881 653 887
rect 595 847 607 881
rect 641 847 653 881
rect 595 841 653 847
rect 787 881 845 887
rect 787 847 799 881
rect 833 847 845 881
rect 787 841 845 847
rect 979 881 1037 887
rect 979 847 991 881
rect 1025 847 1037 881
rect 979 841 1037 847
rect 1171 881 1229 887
rect 1171 847 1183 881
rect 1217 847 1229 881
rect 1171 841 1229 847
rect 1363 881 1421 887
rect 1363 847 1375 881
rect 1409 847 1421 881
rect 1363 841 1421 847
rect -1463 788 -1417 800
rect -1463 -788 -1457 788
rect -1423 -788 -1417 788
rect -1463 -800 -1417 -788
rect -1367 788 -1321 800
rect -1367 -788 -1361 788
rect -1327 -788 -1321 788
rect -1367 -800 -1321 -788
rect -1271 788 -1225 800
rect -1271 -788 -1265 788
rect -1231 -788 -1225 788
rect -1271 -800 -1225 -788
rect -1175 788 -1129 800
rect -1175 -788 -1169 788
rect -1135 -788 -1129 788
rect -1175 -800 -1129 -788
rect -1079 788 -1033 800
rect -1079 -788 -1073 788
rect -1039 -788 -1033 788
rect -1079 -800 -1033 -788
rect -983 788 -937 800
rect -983 -788 -977 788
rect -943 -788 -937 788
rect -983 -800 -937 -788
rect -887 788 -841 800
rect -887 -788 -881 788
rect -847 -788 -841 788
rect -887 -800 -841 -788
rect -791 788 -745 800
rect -791 -788 -785 788
rect -751 -788 -745 788
rect -791 -800 -745 -788
rect -695 788 -649 800
rect -695 -788 -689 788
rect -655 -788 -649 788
rect -695 -800 -649 -788
rect -599 788 -553 800
rect -599 -788 -593 788
rect -559 -788 -553 788
rect -599 -800 -553 -788
rect -503 788 -457 800
rect -503 -788 -497 788
rect -463 -788 -457 788
rect -503 -800 -457 -788
rect -407 788 -361 800
rect -407 -788 -401 788
rect -367 -788 -361 788
rect -407 -800 -361 -788
rect -311 788 -265 800
rect -311 -788 -305 788
rect -271 -788 -265 788
rect -311 -800 -265 -788
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect 265 788 311 800
rect 265 -788 271 788
rect 305 -788 311 788
rect 265 -800 311 -788
rect 361 788 407 800
rect 361 -788 367 788
rect 401 -788 407 788
rect 361 -800 407 -788
rect 457 788 503 800
rect 457 -788 463 788
rect 497 -788 503 788
rect 457 -800 503 -788
rect 553 788 599 800
rect 553 -788 559 788
rect 593 -788 599 788
rect 553 -800 599 -788
rect 649 788 695 800
rect 649 -788 655 788
rect 689 -788 695 788
rect 649 -800 695 -788
rect 745 788 791 800
rect 745 -788 751 788
rect 785 -788 791 788
rect 745 -800 791 -788
rect 841 788 887 800
rect 841 -788 847 788
rect 881 -788 887 788
rect 841 -800 887 -788
rect 937 788 983 800
rect 937 -788 943 788
rect 977 -788 983 788
rect 937 -800 983 -788
rect 1033 788 1079 800
rect 1033 -788 1039 788
rect 1073 -788 1079 788
rect 1033 -800 1079 -788
rect 1129 788 1175 800
rect 1129 -788 1135 788
rect 1169 -788 1175 788
rect 1129 -800 1175 -788
rect 1225 788 1271 800
rect 1225 -788 1231 788
rect 1265 -788 1271 788
rect 1225 -800 1271 -788
rect 1321 788 1367 800
rect 1321 -788 1327 788
rect 1361 -788 1367 788
rect 1321 -800 1367 -788
rect 1417 788 1463 800
rect 1417 -788 1423 788
rect 1457 -788 1463 788
rect 1417 -800 1463 -788
rect -1421 -847 -1363 -841
rect -1421 -881 -1409 -847
rect -1375 -881 -1363 -847
rect -1421 -887 -1363 -881
rect -1229 -847 -1171 -841
rect -1229 -881 -1217 -847
rect -1183 -881 -1171 -847
rect -1229 -887 -1171 -881
rect -1037 -847 -979 -841
rect -1037 -881 -1025 -847
rect -991 -881 -979 -847
rect -1037 -887 -979 -881
rect -845 -847 -787 -841
rect -845 -881 -833 -847
rect -799 -881 -787 -847
rect -845 -887 -787 -881
rect -653 -847 -595 -841
rect -653 -881 -641 -847
rect -607 -881 -595 -847
rect -653 -887 -595 -881
rect -461 -847 -403 -841
rect -461 -881 -449 -847
rect -415 -881 -403 -847
rect -461 -887 -403 -881
rect -269 -847 -211 -841
rect -269 -881 -257 -847
rect -223 -881 -211 -847
rect -269 -887 -211 -881
rect -77 -847 -19 -841
rect -77 -881 -65 -847
rect -31 -881 -19 -847
rect -77 -887 -19 -881
rect 115 -847 173 -841
rect 115 -881 127 -847
rect 161 -881 173 -847
rect 115 -887 173 -881
rect 307 -847 365 -841
rect 307 -881 319 -847
rect 353 -881 365 -847
rect 307 -887 365 -881
rect 499 -847 557 -841
rect 499 -881 511 -847
rect 545 -881 557 -847
rect 499 -887 557 -881
rect 691 -847 749 -841
rect 691 -881 703 -847
rect 737 -881 749 -847
rect 691 -887 749 -881
rect 883 -847 941 -841
rect 883 -881 895 -847
rect 929 -881 941 -847
rect 883 -887 941 -881
rect 1075 -847 1133 -841
rect 1075 -881 1087 -847
rect 1121 -881 1133 -847
rect 1075 -887 1133 -881
rect 1267 -847 1325 -841
rect 1267 -881 1279 -847
rect 1313 -881 1325 -847
rect 1267 -887 1325 -881
<< properties >>
string FIXED_BBOX -1554 -966 1554 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8 l 0.15 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
