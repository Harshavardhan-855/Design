magic
tech sky130A
magscale 1 2
timestamp 1708427080
<< checkpaint >>
rect -1260 1003 1460 1460
rect 3766 1003 7606 1822
rect -1260 -3260 7606 1003
<< error_s >>
rect 8416 8156 8442 8158
rect 8450 8156 8476 8158
rect 11280 8156 11306 8158
rect 11314 8156 11340 8158
rect 7560 8122 12034 8156
rect 7468 8060 7498 8122
rect 7502 8060 7536 8122
rect 7540 8060 7574 8122
rect 7578 8060 7612 8122
rect 7616 8060 7650 8122
rect 7692 8076 7704 8122
rect 7460 8054 7652 8060
rect 7460 8042 7666 8054
rect 7688 8042 7690 8060
rect 7692 8042 7726 8076
rect 7756 8048 7762 8118
rect 7784 8048 7790 8118
rect 8416 8042 8442 8122
rect 8450 8042 8476 8122
rect 9083 8042 9129 8054
rect 9852 8042 9878 8122
rect 9886 8042 9912 8122
rect 10519 8042 10565 8054
rect 11280 8042 11306 8122
rect 11314 8042 11340 8122
rect 11872 8054 11902 8122
rect 11868 8042 11902 8054
rect 7460 8033 9063 8042
rect 9083 8033 10499 8042
rect 10519 8033 11902 8042
rect 11906 8033 11940 8122
rect 11944 8033 11978 8122
rect 7460 8022 11978 8033
rect 7468 7810 7498 8022
rect 7502 8017 7536 8022
rect 7540 8017 7574 8022
rect 7578 8017 7612 8022
rect 7616 8017 11978 8022
rect 7502 8008 11978 8017
rect 7502 7999 7828 8008
rect 8847 7999 9075 8008
rect 9083 8002 9300 8008
rect 9852 8006 9878 8008
rect 9886 8006 9912 8008
rect 9083 7999 9264 8002
rect 10283 7999 10511 8008
rect 10519 8002 10738 8008
rect 10519 7999 10700 8002
rect 7502 7996 7844 7999
rect 8847 7996 9280 7999
rect 10283 7996 10716 7999
rect 7502 7983 7828 7996
rect 8847 7983 9272 7996
rect 10283 7983 10710 7996
rect 11719 7983 11978 8008
rect 7502 7810 7536 7983
rect 7540 7949 7762 7983
rect 7540 7810 7574 7949
rect 7578 7810 7612 7949
rect 7616 7936 7676 7949
rect 7680 7936 7752 7949
rect 7756 7936 7762 7949
rect 7784 7936 7790 7983
rect 7794 7936 7828 7983
rect 8888 7974 8966 7983
rect 8888 7937 8890 7958
rect 8894 7936 8928 7974
rect 8932 7936 8966 7974
rect 8970 7949 9112 7983
rect 9116 7949 9188 7983
rect 9216 7974 9272 7983
rect 10320 7974 10402 7983
rect 8970 7936 9188 7949
rect 9230 7936 9264 7974
rect 10330 7936 10364 7974
rect 10368 7936 10402 7974
rect 10406 7949 10548 7983
rect 10552 7949 10624 7983
rect 10650 7974 10710 7983
rect 10406 7936 10624 7949
rect 10666 7936 10700 7974
rect 11766 7936 11800 7983
rect 11804 7936 11838 7983
rect 11842 7936 11978 7983
rect 7616 7933 7768 7936
rect 7778 7933 7844 7936
rect 8878 7933 9204 7936
rect 9214 7933 9280 7936
rect 10314 7933 10640 7936
rect 10650 7933 10716 7936
rect 11750 7933 11978 7936
rect 7616 7924 7666 7933
rect 7692 7924 7726 7933
rect 7756 7930 7762 7933
rect 7784 7930 7790 7933
rect 9060 7930 9129 7933
rect 8860 7924 8890 7930
rect 9055 7924 9075 7930
rect 9083 7924 9129 7930
rect 10496 7926 10511 7933
rect 10491 7924 10511 7926
rect 10519 7924 10565 7933
rect 11868 7924 11902 7933
rect 11906 7924 11940 7933
rect 11944 7924 11978 7933
rect 7616 7899 11978 7924
rect 7616 7890 9063 7899
rect 9083 7892 10511 7899
rect 10519 7892 11902 7899
rect 9083 7890 10512 7892
rect 7616 7878 7666 7890
rect 7692 7878 7726 7890
rect 8854 7884 8864 7890
rect 8892 7884 8902 7890
rect 8930 7884 8940 7890
rect 8968 7884 8978 7890
rect 9006 7884 9054 7890
rect 9083 7884 9129 7890
rect 9142 7884 9152 7890
rect 9180 7884 9190 7890
rect 9218 7884 9228 7890
rect 9256 7884 9304 7890
rect 10284 7884 10286 7890
rect 10322 7884 10324 7890
rect 10360 7884 10362 7890
rect 10398 7884 10400 7890
rect 10436 7884 10476 7890
rect 8836 7882 8854 7884
rect 8864 7882 8892 7884
rect 8902 7882 8930 7884
rect 8940 7882 8968 7884
rect 8978 7882 8996 7884
rect 9083 7882 9142 7884
rect 9152 7882 9180 7884
rect 9190 7882 9218 7884
rect 9228 7882 9246 7884
rect 7616 7810 7650 7878
rect 7692 7810 7704 7878
rect 8854 7856 8864 7882
rect 8892 7856 8902 7882
rect 8930 7856 8940 7882
rect 8968 7856 8978 7882
rect 9006 7856 9054 7882
rect 9083 7878 9129 7882
rect 9104 7856 9114 7878
rect 9142 7856 9152 7882
rect 9180 7856 9190 7882
rect 9218 7856 9228 7882
rect 9256 7856 9304 7882
rect 10258 7862 10284 7884
rect 10286 7862 10322 7884
rect 10324 7862 10360 7884
rect 10362 7862 10398 7884
rect 10400 7862 10426 7884
rect 10490 7862 10512 7890
rect 10518 7890 11902 7892
rect 10518 7884 10565 7890
rect 10592 7884 10594 7890
rect 10630 7884 10632 7890
rect 10668 7884 10670 7890
rect 10706 7884 10746 7890
rect 10518 7878 10592 7884
rect 10518 7862 10554 7878
rect 10556 7862 10592 7878
rect 10594 7862 10630 7884
rect 10632 7862 10668 7884
rect 10670 7862 10696 7884
rect 10284 7856 10286 7862
rect 10322 7856 10324 7862
rect 10360 7856 10362 7862
rect 10398 7856 10400 7862
rect 10436 7856 10476 7862
rect 10554 7856 10556 7862
rect 10592 7856 10594 7862
rect 10630 7856 10632 7862
rect 10668 7856 10670 7862
rect 10706 7856 10746 7862
rect 11654 7810 11674 7884
rect 11682 7810 11702 7884
rect 11868 7878 11902 7890
rect 11872 7810 11902 7878
rect 11906 7810 11940 7899
rect 11944 7810 11978 7899
rect 11982 7810 12016 8122
rect 12020 7999 12054 8122
rect 12020 7983 12050 7999
rect 12020 7949 12044 7983
rect 12020 7933 12050 7949
rect 12020 7810 12054 7933
rect 12096 7810 12108 8122
rect 7560 7776 12034 7810
rect 7560 7674 8162 7708
rect 7468 7022 7498 7674
rect 7502 7566 7536 7674
rect 7540 7566 7574 7674
rect 7578 7566 7612 7674
rect 7616 7606 7650 7674
rect 7692 7628 7704 7674
rect 7616 7594 7666 7606
rect 7692 7594 7726 7628
rect 7820 7600 7846 7634
rect 7848 7600 7884 7634
rect 7886 7600 7922 7634
rect 7924 7600 7960 7634
rect 7962 7600 7988 7634
rect 8000 7606 8030 7674
rect 7996 7594 8030 7606
rect 7616 7582 8030 7594
rect 8034 7582 8068 7674
rect 8072 7634 8122 7674
rect 8184 7672 11518 7706
rect 8168 7634 8198 7672
rect 8202 7634 8252 7672
rect 8072 7610 8144 7634
rect 8146 7612 8252 7634
rect 8316 7626 8328 7672
rect 8146 7610 8258 7612
rect 8072 7583 8274 7610
rect 8316 7592 8350 7626
rect 9824 7604 9854 7672
rect 9820 7592 9854 7604
rect 8283 7583 9854 7592
rect 9858 7583 9892 7672
rect 9896 7583 9930 7672
rect 8072 7582 9930 7583
rect 7616 7566 9930 7582
rect 7502 7558 9930 7566
rect 7502 7554 8492 7558
rect 7502 7550 7846 7554
rect 7847 7552 8492 7554
rect 7847 7550 8452 7552
rect 7502 7544 7828 7550
rect 7847 7549 8464 7550
rect 7847 7546 8468 7549
rect 7502 7532 7834 7544
rect 7847 7533 8464 7546
rect 9671 7533 9930 7558
rect 9934 7567 9968 7672
rect 9972 7604 10006 7672
rect 10048 7626 10060 7672
rect 9972 7592 10022 7604
rect 10048 7592 10082 7626
rect 11356 7604 11386 7672
rect 11352 7592 11386 7604
rect 9972 7583 11386 7592
rect 11390 7583 11424 7672
rect 11428 7598 11462 7672
rect 11426 7583 11462 7598
rect 9972 7578 11462 7583
rect 11466 7578 11500 7672
rect 9972 7567 11500 7578
rect 9934 7558 11500 7567
rect 9934 7552 10220 7558
rect 9934 7549 10184 7552
rect 9934 7546 10200 7549
rect 9934 7533 10192 7546
rect 11203 7533 11500 7558
rect 7847 7532 8388 7533
rect 7502 7022 7536 7532
rect 7540 7170 7760 7532
rect 7788 7522 7834 7532
rect 7888 7522 8388 7532
rect 7794 7170 7828 7522
rect 7894 7170 7928 7522
rect 7932 7170 7966 7522
rect 7970 7499 8388 7522
rect 7970 7482 8198 7499
rect 8202 7486 8388 7499
rect 8408 7524 8464 7533
rect 9712 7524 10192 7533
rect 11242 7524 11500 7533
rect 8408 7508 8416 7524
rect 8418 7508 8452 7524
rect 9718 7508 9752 7524
rect 9756 7508 9790 7524
rect 9794 7508 10116 7524
rect 10150 7508 10184 7524
rect 11250 7508 11284 7524
rect 11288 7508 11322 7524
rect 11326 7508 11500 7524
rect 8408 7486 8464 7508
rect 9712 7499 10116 7508
rect 9712 7486 9930 7499
rect 8202 7483 8392 7486
rect 8402 7483 8468 7486
rect 9702 7483 9930 7486
rect 8202 7482 8274 7483
rect 8296 7482 8388 7483
rect 8408 7482 8464 7483
rect 7970 7474 8274 7482
rect 8316 7480 8350 7482
rect 9820 7480 9854 7483
rect 8296 7474 8492 7480
rect 9684 7474 9854 7480
rect 9858 7474 9892 7483
rect 9896 7474 9930 7483
rect 7970 7449 9930 7474
rect 7970 7426 8274 7449
rect 8283 7440 9854 7449
rect 7970 7360 8198 7426
rect 8202 7422 8274 7426
rect 8316 7428 8350 7440
rect 8462 7434 8498 7440
rect 9820 7428 9854 7440
rect 8202 7360 8258 7422
rect 8316 7360 8328 7428
rect 8462 7406 8498 7426
rect 9824 7360 9854 7428
rect 9858 7360 9892 7449
rect 9896 7360 9930 7449
rect 9934 7360 9968 7499
rect 9972 7486 10032 7499
rect 10036 7486 10108 7499
rect 10118 7486 10192 7508
rect 11242 7486 11500 7508
rect 9972 7483 10124 7486
rect 10134 7483 10200 7486
rect 11234 7483 11500 7486
rect 9972 7480 10042 7483
rect 10048 7480 10082 7483
rect 11242 7482 11500 7483
rect 11352 7480 11386 7482
rect 11390 7480 11424 7482
rect 11428 7480 11500 7482
rect 9972 7474 10022 7480
rect 10042 7474 10082 7480
rect 10118 7474 10220 7480
rect 11214 7474 11500 7480
rect 9972 7454 11500 7474
rect 9972 7449 11462 7454
rect 9972 7440 11386 7449
rect 9972 7434 10022 7440
rect 9972 7428 10042 7434
rect 9972 7360 10006 7428
rect 10020 7362 10042 7428
rect 10048 7428 10082 7440
rect 10048 7362 10070 7428
rect 10100 7362 10118 7434
rect 10128 7362 10146 7434
rect 10328 7362 10340 7434
rect 10356 7362 10368 7434
rect 11352 7428 11386 7440
rect 10048 7360 10060 7362
rect 11356 7360 11386 7428
rect 11390 7360 11424 7449
rect 11426 7434 11462 7449
rect 11428 7360 11462 7434
rect 11466 7360 11500 7454
rect 11504 7549 11538 7672
rect 11504 7533 11534 7549
rect 11504 7499 11528 7533
rect 11504 7483 11534 7499
rect 11504 7360 11538 7483
rect 11580 7360 11592 7672
rect 7970 7326 8182 7360
rect 8184 7326 11518 7360
rect 7970 7286 8106 7326
rect 8110 7286 8144 7326
rect 8148 7286 8182 7326
rect 8224 7286 8258 7326
rect 7970 7282 8294 7286
rect 7970 7250 8320 7282
rect 7970 7216 9558 7250
rect 7970 7188 8320 7216
rect 7970 7170 8294 7188
rect 7540 7164 7836 7170
rect 7540 7022 7574 7164
rect 7578 7022 7612 7164
rect 7616 7152 7836 7164
rect 7888 7152 8294 7170
rect 7616 7148 7676 7152
rect 7680 7148 7752 7152
rect 7794 7148 7828 7152
rect 7894 7148 7928 7152
rect 7932 7148 7966 7152
rect 7970 7148 8294 7152
rect 8334 7182 8346 7216
rect 8334 7148 8368 7182
rect 9396 7175 9426 7216
rect 9392 7148 9426 7175
rect 7616 7142 7666 7148
rect 7692 7142 7726 7148
rect 7996 7142 8030 7148
rect 7616 7136 8030 7142
rect 8034 7136 8068 7148
rect 8070 7136 9426 7148
rect 7616 7114 9426 7136
rect 7616 7102 8030 7114
rect 7616 7090 7666 7102
rect 7692 7090 7726 7102
rect 7996 7090 8030 7102
rect 7616 7022 7650 7090
rect 7692 7022 7704 7090
rect 8000 7022 8030 7090
rect 8034 7022 8068 7114
rect 8070 7075 8294 7114
rect 8296 7075 8330 7080
rect 8070 7064 8330 7075
rect 8070 7022 8294 7064
rect 7560 6988 8294 7022
rect 8070 6952 8294 6988
rect 8110 6736 8140 6952
rect 8144 6736 8178 6952
rect 8182 6876 8254 6952
rect 8182 6736 8216 6876
rect 8220 6872 8254 6876
rect 8258 6872 8292 6952
rect 8296 6872 8330 7064
rect 8334 7075 8368 7114
rect 8372 7075 8402 7080
rect 9282 7075 9312 7080
rect 9316 7075 9350 7080
rect 9354 7075 9388 7080
rect 8334 7064 8406 7075
rect 8437 7064 8482 7075
rect 9267 7064 9388 7075
rect 8220 6838 8292 6872
rect 8334 6838 8368 7064
rect 8372 6888 8406 7064
rect 8448 6888 8482 7064
rect 9278 6888 9312 7064
rect 8372 6872 8402 6888
rect 9282 6872 9312 6888
rect 9316 6872 9350 7064
rect 9354 6872 9388 7064
rect 9392 6838 9426 7114
rect 8220 6736 8254 6838
rect 8258 6804 9426 6838
rect 8258 6736 8292 6804
rect 8334 6788 8368 6804
rect 8334 6736 8346 6788
rect 8357 6777 8368 6788
rect 9392 6777 9426 6804
rect 9396 6754 9426 6777
rect 9430 6736 9464 7216
rect 9468 7076 9502 7216
rect 9506 7098 9540 7216
rect 9506 7076 9536 7098
rect 9544 7076 9578 7216
rect 9620 7154 9632 7216
rect 9620 7098 9654 7154
rect 10328 7098 10340 7306
rect 10356 7098 10368 7306
rect 9468 7064 9578 7076
rect 9586 7064 11538 7098
rect 9468 6959 9600 7064
rect 9604 7002 9654 7064
rect 9718 7018 9730 7064
rect 9718 7002 9752 7018
rect 9604 6984 9676 7002
rect 9718 6996 9730 7002
rect 9948 6996 9978 7064
rect 9718 6984 9752 6996
rect 9944 6984 9978 6996
rect 9604 6975 9978 6984
rect 9982 6975 10016 7064
rect 10020 6975 10054 7064
rect 9604 6959 10054 6975
rect 9468 6950 10054 6959
rect 9468 6941 9778 6950
rect 9782 6941 10054 6950
rect 9468 6938 10054 6941
rect 9468 6925 9778 6938
rect 9782 6925 10054 6938
rect 10058 6959 10092 7064
rect 10096 6996 10130 7064
rect 10172 7018 10184 7064
rect 10172 7002 10206 7018
rect 10172 6996 10184 7002
rect 10096 6984 10146 6996
rect 10172 6984 10206 6996
rect 10328 6990 10340 7064
rect 10356 6990 10368 7064
rect 10662 6996 10692 7064
rect 10658 6984 10692 6996
rect 10096 6975 10692 6984
rect 10696 6975 10730 7064
rect 10734 6975 10768 7064
rect 10096 6959 10768 6975
rect 10058 6950 10768 6959
rect 10058 6941 10232 6950
rect 10236 6941 10308 6950
rect 10058 6938 10324 6941
rect 10058 6925 10232 6938
rect 10236 6925 10308 6938
rect 10518 6925 10768 6950
rect 10772 6959 10806 7064
rect 10810 6996 10844 7064
rect 10886 7018 10898 7064
rect 10886 7002 10920 7018
rect 10886 6996 10898 7002
rect 11376 6996 11406 7064
rect 10810 6984 10860 6996
rect 10886 6984 10920 6996
rect 11372 6984 11406 6996
rect 10810 6975 11406 6984
rect 11410 6975 11444 7064
rect 11448 7022 11482 7064
rect 11486 7022 11520 7064
rect 11446 6975 11520 7022
rect 10810 6959 11520 6975
rect 10772 6950 11520 6959
rect 10772 6941 10946 6950
rect 10950 6941 11022 6950
rect 11232 6946 11520 6950
rect 10772 6938 11038 6941
rect 10772 6925 10946 6938
rect 10950 6925 11022 6938
rect 11232 6925 11482 6946
rect 9468 6891 9788 6925
rect 9468 6814 9600 6891
rect 9468 6798 9502 6814
rect 9506 6798 9540 6814
rect 9544 6798 9600 6814
rect 9468 6788 9498 6798
rect 9468 6736 9518 6788
rect 9570 6754 9600 6798
rect 9604 6878 9702 6891
rect 9706 6878 9778 6891
rect 9784 6878 9788 6891
rect 9812 6878 9816 6925
rect 9820 6878 9876 6925
rect 9880 6878 9914 6925
rect 9918 6891 10240 6925
rect 9918 6878 10054 6891
rect 9604 6875 9794 6878
rect 9804 6875 10054 6878
rect 9604 6866 9676 6875
rect 9718 6866 9752 6875
rect 9784 6872 9788 6875
rect 9812 6872 9816 6875
rect 9944 6866 9978 6875
rect 9982 6872 10016 6875
rect 10020 6872 10054 6875
rect 10058 6872 10092 6891
rect 9982 6870 10092 6872
rect 9982 6866 10054 6870
rect 9604 6841 10054 6866
rect 9604 6832 9978 6841
rect 9604 6814 9676 6832
rect 9718 6820 9752 6832
rect 9604 6752 9654 6814
rect 9718 6752 9730 6820
rect 9904 6752 9908 6832
rect 9938 6752 9942 6832
rect 9944 6820 9978 6832
rect 9982 6752 10016 6841
rect 10020 6752 10054 6841
rect 10058 6752 10092 6870
rect 10096 6878 10156 6891
rect 10160 6878 10232 6891
rect 10274 6878 10308 6925
rect 10556 6878 10590 6925
rect 10594 6878 10628 6925
rect 10632 6891 10954 6925
rect 10632 6878 10768 6891
rect 10096 6875 10248 6878
rect 10258 6875 10324 6878
rect 10540 6875 10768 6878
rect 10096 6866 10146 6875
rect 10172 6866 10206 6875
rect 10658 6866 10692 6875
rect 10696 6866 10730 6875
rect 10734 6866 10768 6875
rect 10096 6841 10768 6866
rect 10096 6832 10692 6841
rect 10096 6820 10146 6832
rect 10172 6820 10206 6832
rect 10096 6752 10130 6820
rect 10172 6752 10184 6820
rect 10486 6752 10490 6832
rect 10520 6752 10524 6832
rect 10658 6820 10692 6832
rect 10662 6752 10692 6820
rect 10696 6752 10730 6841
rect 10734 6752 10768 6841
rect 10772 6752 10806 6891
rect 10810 6878 10870 6891
rect 10874 6878 10946 6891
rect 10988 6878 11022 6925
rect 11270 6878 11304 6925
rect 11308 6878 11342 6925
rect 11346 6878 11482 6925
rect 10810 6875 10962 6878
rect 10972 6875 11038 6878
rect 11254 6875 11482 6878
rect 10810 6866 10860 6875
rect 10886 6866 10920 6875
rect 11372 6866 11406 6875
rect 11410 6866 11444 6875
rect 11448 6866 11482 6875
rect 10810 6841 11482 6866
rect 10810 6832 11406 6841
rect 10810 6820 10860 6832
rect 10886 6820 10920 6832
rect 10810 6752 10844 6820
rect 10886 6752 10898 6820
rect 11208 6752 11212 6832
rect 11242 6752 11246 6832
rect 11372 6820 11406 6832
rect 11376 6754 11406 6820
rect 11410 6754 11444 6841
rect 11448 6754 11482 6841
rect 11486 6754 11520 6946
rect 11524 6941 11558 7064
rect 11524 6925 11554 6941
rect 11524 6891 11548 6925
rect 11524 6875 11554 6891
rect 11524 6754 11558 6875
rect 11364 6752 11558 6754
rect 8202 6702 9558 6736
rect 9586 6718 11558 6752
rect 11592 6718 11596 6754
rect 11600 6752 11612 7064
rect 11654 7054 11674 7776
rect 11682 7054 11702 7776
rect 11796 7182 12118 7306
rect 9904 6716 9908 6718
rect 9938 6716 9942 6718
rect 10486 6714 10490 6718
rect 10520 6714 10524 6718
rect 2191 3481 2457 3483
rect 2571 3475 2664 3483
rect 1777 3452 1862 3453
rect 1408 3415 1423 3449
rect 1462 3434 1515 3449
rect 1558 3447 1573 3449
rect 1446 3425 1515 3434
rect 1554 3431 1595 3447
rect 1767 3436 1862 3452
rect 1949 3449 2053 3453
rect 1446 3405 1512 3425
rect 1554 3415 1607 3431
rect 1524 3405 1529 3415
rect 1554 3406 1599 3415
rect 1370 3346 1372 3384
rect 1398 3374 1400 3384
rect 1446 3382 1496 3405
rect 1412 3348 1429 3381
rect 1454 3371 1463 3382
rect 1523 3379 1553 3405
rect 1554 3396 1595 3406
rect 1469 3375 1523 3379
rect 1420 3305 1429 3348
rect 1482 3364 1523 3375
rect 1482 3352 1512 3364
rect 1454 3333 1463 3337
rect 1482 3333 1523 3352
rect 1524 3337 1529 3379
rect 1558 3375 1563 3396
rect 1597 3379 1604 3406
rect 1584 3375 1605 3379
rect 1631 3375 1638 3378
rect 1685 3375 1696 3378
rect 1719 3375 1730 3412
rect 1558 3337 1749 3375
rect 1561 3333 1749 3337
rect 1780 3333 1811 3415
rect 1854 3385 1862 3436
rect 1925 3425 2053 3449
rect 2079 3425 2087 3453
rect 2590 3449 2623 3453
rect 2159 3447 2457 3449
rect 2571 3441 2711 3449
rect 1873 3385 1879 3415
rect 1925 3411 1980 3425
rect 2415 3415 2423 3427
rect 2590 3425 2623 3441
rect 2642 3431 2653 3441
rect 2677 3431 2711 3441
rect 2603 3415 2623 3425
rect 1884 3395 1912 3411
rect 1925 3397 1959 3411
rect 1949 3395 1954 3397
rect 1926 3385 1954 3395
rect 1981 3385 2011 3411
rect 2124 3397 2156 3413
rect 2158 3397 2190 3413
rect 2241 3399 2248 3411
rect 2241 3397 2375 3399
rect 1839 3381 1882 3385
rect 1814 3370 1882 3381
rect 1889 3383 2051 3385
rect 2072 3383 2119 3385
rect 1889 3379 2119 3383
rect 1814 3333 1845 3370
rect 1854 3333 1882 3370
rect 1907 3373 2119 3379
rect 1907 3370 2017 3373
rect 1907 3363 1913 3370
rect 1926 3363 2017 3370
rect 2022 3363 2119 3373
rect 1907 3349 2119 3363
rect 1907 3333 2121 3349
rect 2122 3333 2156 3397
rect 2157 3388 2375 3397
rect 2415 3393 2425 3415
rect 2423 3388 2425 3393
rect 2457 3388 2459 3415
rect 2611 3413 2623 3415
rect 2641 3415 2711 3431
rect 2760 3415 2790 3453
rect 3500 3449 3520 3496
rect 3554 3465 3588 3496
rect 3534 3460 3568 3462
rect 3534 3449 3622 3460
rect 2798 3415 2855 3439
rect 2857 3415 2895 3449
rect 3106 3415 3143 3441
rect 3240 3415 3263 3449
rect 3296 3430 3355 3449
rect 3278 3415 3355 3430
rect 2641 3411 2677 3415
rect 2714 3411 2743 3415
rect 2641 3397 2675 3411
rect 2684 3388 2743 3411
rect 2748 3411 2790 3415
rect 2748 3388 2777 3411
rect 2792 3405 2822 3411
rect 2798 3388 2821 3405
rect 2857 3392 2891 3415
rect 2965 3397 2971 3415
rect 2157 3385 2845 3388
rect 2857 3385 2900 3392
rect 2903 3385 2991 3397
rect 2157 3384 2991 3385
rect 2158 3369 2190 3384
rect 2196 3370 2218 3384
rect 2268 3375 2300 3384
rect 2363 3377 2415 3384
rect 2423 3377 2425 3384
rect 2457 3377 2459 3384
rect 2490 3383 2556 3384
rect 2490 3377 2581 3383
rect 2339 3375 2581 3377
rect 2211 3369 2218 3370
rect 2245 3369 2581 3375
rect 2158 3367 2581 3369
rect 2158 3363 2525 3367
rect 2537 3363 2581 3367
rect 2630 3381 2743 3384
rect 2630 3370 2684 3381
rect 2630 3365 2677 3370
rect 2714 3369 2743 3381
rect 2745 3383 2963 3384
rect 2745 3373 2889 3383
rect 2748 3370 2889 3373
rect 2748 3369 2858 3370
rect 2630 3363 2653 3365
rect 2714 3363 2858 3369
rect 2863 3369 2889 3370
rect 2891 3375 2932 3383
rect 2944 3375 2963 3383
rect 2965 3375 2971 3384
rect 2999 3375 3005 3415
rect 3068 3391 3143 3415
rect 3106 3385 3143 3391
rect 3166 3385 3174 3415
rect 3200 3385 3208 3415
rect 3278 3388 3330 3415
rect 3335 3385 3350 3415
rect 2891 3370 3019 3375
rect 2891 3369 2917 3370
rect 2921 3369 3019 3370
rect 2863 3367 2876 3369
rect 2158 3360 2669 3363
rect 2714 3360 2866 3363
rect 2158 3356 2866 3360
rect 2158 3339 2190 3356
rect 2211 3343 2218 3356
rect 2245 3349 2669 3356
rect 2714 3355 2866 3356
rect 2197 3339 2231 3343
rect 2245 3339 2684 3349
rect 2158 3333 2684 3339
rect 2714 3339 2792 3355
rect 2798 3349 2821 3355
rect 2832 3349 2866 3355
rect 2868 3349 2876 3367
rect 2902 3361 3019 3369
rect 2902 3356 3043 3361
rect 3068 3357 3072 3381
rect 3106 3379 3174 3385
rect 3198 3379 3260 3385
rect 3290 3379 3350 3385
rect 3369 3379 3384 3415
rect 3408 3407 3416 3441
rect 3520 3431 3622 3449
rect 3402 3391 3416 3407
rect 3428 3391 3452 3425
rect 3408 3385 3416 3391
rect 3393 3379 3434 3385
rect 3444 3379 3452 3391
rect 3466 3385 3664 3421
rect 3458 3379 3664 3385
rect 3106 3378 3664 3379
rect 3106 3377 3804 3378
rect 3101 3375 3804 3377
rect 3101 3362 3106 3375
rect 2714 3333 2832 3339
rect 2868 3333 2883 3349
rect 2902 3343 2917 3356
rect 2921 3343 3043 3356
rect 2902 3339 3043 3343
rect 2917 3333 3043 3339
rect 3069 3333 3072 3357
rect 3103 3333 3106 3353
rect 3147 3333 3804 3375
rect 1387 3271 1431 3289
rect 1378 3266 1431 3271
rect 1437 3266 3804 3333
rect 1378 3247 3804 3266
rect 1408 3240 3804 3247
rect 1344 3213 1391 3237
rect 1437 3235 3804 3240
rect 1431 3206 3804 3235
rect 1431 3184 1436 3206
rect 1437 3197 3804 3206
rect 1447 3184 1553 3197
rect 1608 3193 1644 3197
rect 1700 3195 1776 3197
rect 1782 3195 1820 3197
rect 1700 3193 1820 3195
rect 1975 3193 2039 3197
rect 2121 3193 2176 3197
rect 2218 3193 2248 3197
rect 2325 3193 2328 3197
rect 2339 3193 2377 3197
rect 2387 3193 2449 3197
rect 2514 3193 2544 3197
rect 2646 3193 2676 3197
rect 2680 3193 2714 3197
rect 2743 3193 2760 3197
rect 2777 3193 2822 3197
rect 2864 3195 2933 3197
rect 2868 3193 2918 3195
rect 2958 3193 2967 3197
rect 2981 3193 2996 3197
rect 3071 3193 3101 3197
rect 3153 3193 3158 3197
rect 3168 3193 3198 3197
rect 3222 3193 3252 3197
rect 3259 3195 3293 3197
rect 3312 3195 3327 3197
rect 3260 3193 3290 3195
rect 3306 3193 3332 3195
rect 3344 3193 3374 3197
rect 3384 3195 3420 3197
rect 3428 3193 3474 3197
rect 3478 3193 3520 3197
rect 3612 3194 3804 3197
rect 1349 3161 1553 3184
rect 1557 3180 1644 3193
rect 1649 3184 1820 3193
rect 1557 3161 1623 3180
rect 1332 3127 1347 3161
rect 1349 3159 1623 3161
rect 1649 3172 1808 3184
rect 1649 3159 1823 3172
rect 1833 3167 1899 3193
rect 1925 3172 2011 3193
rect 2017 3172 2083 3193
rect 1925 3167 2083 3172
rect 1833 3165 2083 3167
rect 2109 3177 2176 3193
rect 2109 3172 2175 3177
rect 2109 3165 2180 3172
rect 2201 3165 2267 3193
rect 1833 3159 2267 3165
rect 2293 3186 2377 3193
rect 2385 3186 2451 3193
rect 2293 3159 2451 3186
rect 2477 3174 2544 3193
rect 2569 3174 2635 3193
rect 2477 3165 2638 3174
rect 2661 3172 2727 3193
rect 2753 3176 2822 3193
rect 2828 3184 3003 3193
rect 3029 3184 3101 3193
rect 3121 3184 3198 3193
rect 2828 3176 3198 3184
rect 2661 3165 2729 3172
rect 1349 3152 1559 3159
rect 1349 3145 1473 3152
rect 1478 3145 1559 3152
rect 1349 3127 1559 3145
rect 1589 3127 1623 3159
rect 1681 3157 1823 3159
rect 1844 3157 2026 3159
rect 1681 3148 1807 3157
rect 1681 3127 1715 3148
rect 1752 3127 1807 3148
rect 1844 3137 1991 3157
rect 2003 3137 2011 3157
rect 1844 3135 1904 3137
rect 1844 3127 1937 3135
rect 1943 3127 1991 3137
rect 2049 3127 2113 3159
rect 2120 3157 2267 3159
rect 1340 3122 1559 3127
rect 1563 3122 1593 3127
rect 1340 3109 1593 3122
rect 1752 3111 1786 3127
rect 1797 3111 1810 3127
rect 1837 3123 1937 3127
rect 1837 3119 1883 3123
rect 1340 3107 1485 3109
rect 1515 3107 1593 3109
rect 1340 3103 1420 3107
rect 1370 3094 1420 3103
rect 1306 3069 1353 3093
rect 1378 3083 1387 3094
rect 1447 3091 1477 3107
rect 1485 3091 1515 3107
rect 1523 3091 1559 3107
rect 1393 3076 1447 3091
rect 1477 3090 1559 3091
rect 1563 3090 1593 3107
rect 1735 3097 1803 3111
rect 1837 3109 1844 3119
rect 1849 3109 1883 3119
rect 1837 3097 1878 3109
rect 1903 3101 1937 3123
rect 1905 3097 1937 3101
rect 1941 3097 1973 3127
rect 1975 3097 2005 3127
rect 2009 3125 2039 3127
rect 2083 3117 2113 3127
rect 2135 3127 2175 3157
rect 2135 3125 2155 3127
rect 2180 3125 2210 3157
rect 2218 3127 2267 3157
rect 2218 3125 2248 3127
rect 2135 3117 2254 3125
rect 2275 3121 2288 3125
rect 2048 3109 2080 3117
rect 2082 3109 2114 3117
rect 2135 3109 2155 3117
rect 2180 3111 2210 3117
rect 2218 3111 2248 3117
rect 2275 3111 2289 3121
rect 2325 3111 2394 3159
rect 2417 3138 2451 3159
rect 2476 3157 2638 3165
rect 2646 3157 2729 3165
rect 2753 3161 3198 3176
rect 2753 3159 2925 3161
rect 2937 3159 3198 3161
rect 3213 3161 3293 3193
rect 3305 3184 3374 3193
rect 3397 3187 3463 3193
rect 3390 3185 3463 3187
rect 3213 3159 3290 3161
rect 2754 3157 2925 3159
rect 2417 3127 2461 3138
rect 2415 3126 2461 3127
rect 2169 3109 2299 3111
rect 2046 3097 2080 3109
rect 2081 3100 2299 3109
rect 2325 3105 2411 3111
rect 2325 3100 2377 3105
rect 2381 3100 2411 3105
rect 2414 3100 2461 3126
rect 2476 3100 2506 3157
rect 2509 3127 2561 3157
rect 2566 3143 2592 3157
rect 2601 3143 2635 3157
rect 2565 3127 2635 3143
rect 2516 3123 2608 3127
rect 2633 3123 2642 3127
rect 2516 3109 2642 3123
rect 2516 3101 2592 3109
rect 2516 3100 2548 3101
rect 2557 3100 2592 3101
rect 2599 3100 2642 3109
rect 2646 3100 2676 3157
rect 2684 3151 2727 3157
rect 2754 3151 2822 3157
rect 2684 3145 2822 3151
rect 2838 3145 2864 3157
rect 2877 3151 2911 3157
rect 2969 3153 3121 3159
rect 3153 3153 3198 3159
rect 3220 3153 3290 3159
rect 2684 3127 2826 3145
rect 2877 3127 2913 3151
rect 2969 3137 3130 3153
rect 2969 3127 3033 3137
rect 2684 3117 2714 3127
rect 2716 3117 2746 3123
rect 2684 3100 2718 3117
rect 2722 3100 2745 3117
rect 2754 3109 2831 3127
rect 2883 3109 2913 3127
rect 2754 3100 2915 3109
rect 2081 3097 2915 3100
rect 1477 3087 1529 3090
rect 1662 3087 1670 3097
rect 1735 3093 1806 3097
rect 1836 3093 2043 3097
rect 1477 3085 1673 3087
rect 1477 3076 1677 3085
rect 1744 3082 1806 3093
rect 1336 3060 1387 3069
rect 1344 3049 1387 3060
rect 1393 3064 1436 3076
rect 1485 3070 1677 3076
rect 1752 3070 1806 3082
rect 1393 3062 1447 3064
rect 1393 3045 1398 3062
rect 1406 3055 1447 3062
rect 1485 3055 1714 3070
rect 1406 3051 1714 3055
rect 1744 3051 1806 3070
rect 1406 3045 1806 3051
rect 1831 3082 2043 3093
rect 1831 3075 1941 3082
rect 1943 3075 2043 3082
rect 1831 3065 2043 3075
rect 1831 3055 1837 3065
rect 1850 3061 2043 3065
rect 2046 3096 2915 3097
rect 2046 3091 2224 3096
rect 2256 3091 2261 3093
rect 2275 3091 2339 3096
rect 2046 3089 2339 3091
rect 2347 3089 2411 3096
rect 2414 3095 2895 3096
rect 2414 3093 2529 3095
rect 2554 3093 2895 3095
rect 2414 3089 2521 3093
rect 2046 3084 2521 3089
rect 2046 3083 2514 3084
rect 1850 3057 2045 3061
rect 1850 3055 1904 3057
rect 1831 3045 1904 3055
rect 1931 3045 2045 3057
rect 2046 3049 2069 3083
rect 2075 3082 2514 3083
rect 2554 3082 2826 3093
rect 2083 3079 2506 3082
rect 2083 3075 2449 3079
rect 2461 3075 2506 3079
rect 2554 3075 2639 3082
rect 2646 3081 2676 3082
rect 2684 3081 2826 3082
rect 2830 3087 2895 3093
rect 2920 3087 2929 3127
rect 2981 3105 3033 3127
rect 3040 3117 3130 3137
rect 3153 3127 3290 3153
rect 3295 3153 3374 3184
rect 3397 3159 3463 3185
rect 3489 3159 3501 3193
rect 3505 3185 3520 3193
rect 3610 3184 3804 3194
rect 3610 3168 3802 3184
rect 3588 3160 3802 3168
rect 3428 3153 3463 3159
rect 3295 3137 3390 3153
rect 3160 3123 3290 3127
rect 3293 3123 3323 3127
rect 3040 3105 3154 3117
rect 2992 3103 3067 3105
rect 3030 3097 3067 3103
rect 3080 3097 3154 3105
rect 2830 3081 2943 3087
rect 2083 3072 2506 3075
rect 2509 3072 2602 3075
rect 2643 3072 2826 3081
rect 2083 3068 2826 3072
rect 2827 3073 2943 3081
rect 2827 3068 2967 3073
rect 2992 3069 2996 3093
rect 3030 3091 3120 3097
rect 3122 3091 3154 3097
rect 3160 3100 3323 3123
rect 3160 3097 3222 3100
rect 3160 3091 3184 3097
rect 3214 3095 3222 3097
rect 3252 3097 3323 3100
rect 3336 3119 3390 3137
rect 3420 3127 3463 3153
rect 3588 3134 3766 3160
rect 3420 3119 3458 3127
rect 3336 3108 3458 3119
rect 3336 3103 3474 3108
rect 3336 3097 3390 3103
rect 3252 3095 3289 3097
rect 3214 3093 3289 3095
rect 3192 3091 3289 3093
rect 3293 3095 3352 3097
rect 3382 3095 3390 3097
rect 3420 3095 3474 3103
rect 3293 3091 3390 3095
rect 3392 3091 3474 3095
rect 3482 3091 3588 3133
rect 3612 3128 3766 3134
rect 3635 3124 3665 3128
rect 3669 3124 3703 3128
rect 3626 3100 3631 3124
rect 3030 3090 3588 3091
rect 3734 3090 3766 3128
rect 3030 3089 3766 3090
rect 3025 3087 3766 3089
rect 3025 3074 3030 3087
rect 2083 3055 2142 3068
rect 2169 3067 2602 3068
rect 2083 3051 2155 3055
rect 2169 3051 2506 3067
rect 2509 3059 2602 3067
rect 2643 3067 2826 3068
rect 2643 3059 2716 3067
rect 2747 3061 2826 3067
rect 2754 3059 2784 3061
rect 2509 3051 2608 3059
rect 2080 3049 2608 3051
rect 2046 3045 2080 3049
rect 2082 3045 2608 3049
rect 2643 3045 2784 3059
rect 2792 3059 2800 3061
rect 2830 3059 2967 3068
rect 2792 3045 2807 3059
rect 2826 3051 2967 3059
rect 2830 3045 2967 3051
rect 2993 3045 2996 3069
rect 3027 3045 3030 3065
rect 3033 3045 3063 3087
rect 3071 3045 3766 3087
rect 1361 3040 3766 3045
rect 1294 2983 1309 3017
rect 1311 3016 3764 3040
rect 1311 2983 3728 3016
rect 1302 2978 3728 2983
rect 1302 2959 3734 2978
rect 12966 2962 13080 2964
rect 1332 2950 3734 2959
rect 1268 2932 1315 2949
rect 1340 2939 1349 2950
rect 1361 2947 3734 2950
rect 1355 2932 3734 2947
rect 1268 2925 3734 2932
rect 12251 2927 12285 2961
rect 12289 2927 12323 2961
rect 12327 2927 12729 2961
rect 12733 2934 12805 2961
rect 12733 2927 12810 2934
rect 1294 2918 3734 2925
rect 1294 2916 1360 2918
rect 1306 2905 1349 2916
rect 1355 2904 1360 2916
rect 1361 2909 3734 2918
rect 1294 2901 1360 2904
rect 1368 2907 1676 2909
rect 1706 2907 1768 2909
rect 1368 2905 1768 2907
rect 1793 2905 1799 2909
rect 1812 2905 1866 2909
rect 1893 2905 2007 2909
rect 2008 2905 2031 2909
rect 2045 2905 2117 2909
rect 1368 2901 2007 2905
rect 2033 2901 2117 2905
rect 2125 2906 2483 2909
rect 2486 2906 2539 2909
rect 2125 2905 2539 2906
rect 2570 2905 2600 2909
rect 2605 2907 2705 2909
rect 2605 2905 2638 2907
rect 2661 2905 2705 2907
rect 2716 2905 2746 2909
rect 2125 2901 2559 2905
rect 2570 2901 2651 2905
rect 2661 2901 2746 2905
rect 2754 2901 2929 2909
rect 2955 2905 2958 2909
rect 2989 2905 2992 2909
rect 2995 2905 3025 2909
rect 2953 2901 3025 2905
rect 3033 2901 3734 2909
rect 1294 2896 3734 2901
rect 1273 2895 3734 2896
rect 1256 2848 1271 2873
rect 1273 2848 3756 2895
rect 12311 2885 12341 2895
rect 12349 2885 12379 2923
rect 12387 2895 12421 2923
rect 12439 2895 12469 2927
rect 12473 2895 12503 2927
rect 12515 2895 12545 2927
rect 12549 2895 12583 2927
rect 12587 2895 12617 2927
rect 12677 2895 12711 2923
rect 12765 2895 12797 2927
rect 12799 2897 12831 2927
rect 12833 2905 12837 2939
rect 12871 2905 12927 2939
rect 12993 2905 13000 2930
rect 13027 2905 13054 2939
rect 12837 2897 12873 2905
rect 12799 2895 12873 2897
rect 12387 2885 12669 2895
rect 12677 2885 12745 2895
rect 12765 2885 12873 2895
rect 12305 2851 12341 2885
rect 12343 2880 12873 2885
rect 12343 2851 12833 2880
rect 1256 2842 3756 2848
rect 1256 2840 3736 2842
rect 1256 2839 3696 2840
rect 1264 2815 3696 2839
rect 3727 2816 3736 2840
rect 12311 2817 12341 2827
rect 12349 2817 12379 2851
rect 12387 2827 12421 2851
rect 12677 2835 12711 2851
rect 12387 2817 12669 2827
rect 12677 2817 12721 2835
rect 1266 2805 3696 2815
rect 1230 2798 3696 2805
rect 1230 2784 1294 2798
rect 1302 2795 1311 2798
rect 1317 2784 3696 2798
rect 1230 2781 1277 2784
rect 1294 2781 3696 2784
rect 12305 2783 12341 2817
rect 12343 2783 12721 2817
rect 1260 2772 3696 2781
rect 1268 2770 3696 2772
rect 1268 2761 1311 2770
rect 1317 2757 1322 2770
rect 1323 2765 3696 2770
rect 1330 2763 1638 2765
rect 1668 2763 1730 2765
rect 1330 2761 1730 2763
rect 1755 2761 1761 2765
rect 1774 2761 1828 2765
rect 1330 2757 1753 2761
rect 1774 2757 1845 2761
rect 1855 2757 1969 2765
rect 1970 2761 1993 2765
rect 2007 2761 2532 2765
rect 2567 2763 2640 2765
rect 2567 2761 2611 2763
rect 1977 2757 2611 2761
rect 2661 2761 2714 2765
rect 2661 2757 2670 2761
rect 2673 2760 2714 2761
rect 2716 2760 2891 2765
rect 2917 2761 2920 2765
rect 2951 2761 2954 2765
rect 2673 2757 2891 2760
rect 2957 2757 2987 2765
rect 2995 2757 3696 2765
rect 1285 2752 3696 2757
rect 1235 2741 3696 2752
rect 12311 2749 12341 2759
rect 12349 2749 12379 2783
rect 12387 2759 12421 2783
rect 12387 2749 12669 2759
rect 12677 2749 12721 2783
rect 1235 2707 3718 2741
rect 12305 2715 12341 2749
rect 12343 2715 12669 2749
rect 12671 2737 12721 2749
rect 12731 2737 12755 2835
rect 12765 2737 12797 2851
rect 12799 2737 12833 2851
rect 12837 2737 12873 2880
rect 12875 2737 12909 2905
rect 12913 2737 12947 2905
rect 12951 2737 12985 2905
rect 13027 2791 13039 2905
rect 12671 2715 12715 2737
rect 12747 2715 12755 2737
rect 1235 2705 3696 2707
rect 1242 2696 3696 2705
rect 1242 2689 3658 2696
rect 1243 2687 3658 2689
rect 1256 2681 3658 2687
rect 1268 2675 3658 2681
rect 1272 2671 3658 2675
rect 1222 2662 1248 2671
rect 1256 2662 3658 2671
rect 12349 2665 12379 2715
rect 12387 2665 12421 2715
rect 12677 2665 12711 2715
rect 12799 2703 12873 2737
rect 12993 2703 13000 2737
rect 13027 2703 13054 2791
rect 12797 2662 12808 2699
rect 12831 2662 12842 2699
rect 1222 2637 1260 2662
rect 1264 2651 3658 2662
rect 1272 2637 3658 2651
rect 1222 2633 3658 2637
rect 1226 2628 3658 2633
rect 1228 2621 3658 2628
rect 1228 2617 1439 2621
rect 1228 2613 1256 2617
rect 1272 2613 1439 2617
rect 1549 2613 1732 2621
rect 1738 2620 1790 2621
rect 1793 2620 1900 2621
rect 1738 2617 1900 2620
rect 1930 2617 1987 2621
rect 1738 2613 1804 2617
rect 1817 2613 1991 2617
rect 2007 2613 2099 2621
rect 2103 2613 2113 2621
rect 2125 2617 2147 2621
rect 2149 2617 3658 2621
rect 2125 2613 3658 2617
rect 1228 2608 3658 2613
rect 1024 2586 1054 2608
rect 1193 2607 3658 2608
rect 12248 2649 12458 2658
rect 12476 2649 12496 2658
rect 12794 2656 12818 2662
rect 12606 2649 12818 2656
rect 12248 2648 12818 2649
rect 12822 2648 12846 2662
rect 12248 2620 12808 2648
rect 12831 2620 12844 2648
rect 12248 2615 12818 2620
rect 1193 2606 3680 2607
rect 1193 2605 3726 2606
rect 1228 2580 3726 2605
rect 12248 2604 12458 2615
rect 12476 2604 12534 2615
rect 12606 2612 12818 2615
rect 12794 2608 12818 2612
rect 12822 2608 12846 2620
rect 12720 2606 12846 2608
rect 12720 2600 12842 2606
rect 12720 2599 12832 2600
rect 12349 2581 12379 2599
rect 12387 2581 12421 2599
rect 1024 2558 1054 2580
rect 1230 2511 1242 2577
rect 1167 2507 1242 2511
rect 1247 2573 3726 2580
rect 1247 2507 2828 2573
rect 2843 2549 2963 2573
rect 2888 2527 2889 2549
rect 2905 2546 2963 2549
rect 2972 2552 3726 2573
rect 12335 2570 12568 2581
rect 2972 2546 3620 2552
rect 1167 2497 2828 2507
rect 2905 2503 3620 2546
rect 1167 2473 1242 2497
rect 1247 2488 2828 2497
rect 2940 2497 3620 2503
rect 3636 2497 3739 2552
rect 1247 2477 2826 2488
rect 1249 2473 1538 2477
rect 1167 2469 1538 2473
rect 1551 2469 1585 2473
rect 1588 2469 1907 2477
rect 1937 2473 2061 2477
rect 1931 2469 2061 2473
rect 2065 2469 2075 2477
rect 2085 2469 2095 2477
rect 2107 2473 2826 2477
rect 2103 2469 2826 2473
rect 1167 2464 2826 2469
rect 1167 2453 2711 2464
rect 1287 2443 1314 2453
rect 1327 2443 1359 2453
rect 1551 2443 1585 2453
rect 1589 2443 1623 2447
rect 1626 2443 1661 2453
rect 1691 2443 1803 2453
rect 1235 2439 1287 2443
rect 1317 2439 1409 2443
rect 1523 2441 1661 2443
rect 1235 2429 1371 2439
rect 1235 2405 1313 2429
rect 1317 2428 1371 2429
rect 1327 2405 1371 2428
rect 1235 2393 1377 2405
rect 1235 2367 1337 2393
rect 1217 2363 1337 2367
rect 1174 2359 1337 2363
rect 1174 2345 1339 2359
rect 1287 2333 1303 2345
rect 1311 2333 1339 2345
rect 1311 2329 1337 2333
rect 1353 2329 1377 2393
rect 1405 2359 1411 2431
rect 1443 2381 1445 2439
rect 1447 2359 1453 2421
rect 1477 2363 1479 2439
rect 1523 2428 1538 2441
rect 1543 2439 1661 2441
rect 1687 2441 1803 2443
rect 1805 2441 1861 2453
rect 1931 2450 1953 2453
rect 1982 2450 2711 2453
rect 1931 2443 2711 2450
rect 1687 2439 1861 2441
rect 1865 2439 2711 2443
rect 2747 2439 2761 2464
rect 2940 2455 3739 2497
rect 12311 2493 12341 2503
rect 12349 2501 12379 2570
rect 12387 2511 12421 2570
rect 12677 2511 12711 2599
rect 12720 2584 12745 2599
rect 12791 2597 12832 2599
rect 12791 2584 12821 2597
rect 12387 2501 12669 2511
rect 12677 2504 12715 2511
rect 12720 2504 13110 2584
rect 12677 2501 13110 2504
rect 12349 2494 12669 2501
rect 12671 2494 13110 2501
rect 12349 2493 13110 2494
rect 12305 2459 12341 2493
rect 12343 2467 13110 2493
rect 12343 2459 12379 2467
rect 12381 2460 13110 2467
rect 12381 2459 12631 2460
rect 12663 2459 12707 2460
rect 2925 2439 3739 2455
rect 1543 2431 1653 2439
rect 1559 2429 1653 2431
rect 1485 2363 1491 2383
rect 1521 2374 1557 2421
rect 1571 2407 1653 2429
rect 1657 2407 1685 2439
rect 1687 2431 1706 2439
rect 1805 2431 1839 2439
rect 1865 2433 2740 2439
rect 1847 2431 2740 2433
rect 1687 2428 2740 2431
rect 1687 2416 1893 2428
rect 1687 2407 1797 2416
rect 1805 2408 1893 2416
rect 1571 2405 1657 2407
rect 1687 2405 1805 2407
rect 1571 2397 1653 2405
rect 1571 2381 1625 2397
rect 1691 2385 1721 2405
rect 1571 2377 1601 2381
rect 1667 2377 1721 2385
rect 1725 2399 1797 2405
rect 1811 2399 1817 2408
rect 1821 2399 1893 2408
rect 1725 2377 1865 2399
rect 1907 2377 1937 2428
rect 1944 2407 2740 2428
rect 1944 2405 2702 2407
rect 2771 2405 2774 2439
rect 2940 2419 3739 2439
rect 12349 2421 12379 2459
rect 12387 2421 12421 2459
rect 1944 2387 2774 2405
rect 2854 2398 2875 2415
rect 2909 2406 2925 2415
rect 2888 2402 2925 2406
rect 2940 2410 3726 2419
rect 12439 2417 12469 2451
rect 12473 2417 12503 2451
rect 12515 2417 12545 2451
rect 12549 2417 12583 2451
rect 12587 2417 12617 2451
rect 12677 2421 12711 2459
rect 12720 2417 13110 2460
rect 2940 2407 3622 2410
rect 3636 2407 3726 2410
rect 2940 2402 3726 2407
rect 1944 2377 2780 2387
rect 2888 2384 3726 2402
rect 2888 2383 3719 2384
rect 12251 2383 12285 2417
rect 12289 2383 12323 2417
rect 12327 2383 13110 2417
rect 2888 2381 3688 2383
rect 1571 2374 2780 2377
rect 1521 2373 2780 2374
rect 1521 2367 2665 2373
rect 2670 2367 2780 2373
rect 2902 2379 3688 2381
rect 2902 2372 3582 2379
rect 1521 2363 2780 2367
rect 2888 2363 3582 2372
rect 1387 2329 1411 2359
rect 1477 2333 1517 2363
rect 1521 2359 3582 2363
rect 1583 2333 1623 2359
rect 1626 2333 1643 2359
rect 1667 2355 1698 2359
rect 1725 2355 1831 2359
rect 1667 2333 1697 2355
rect 1721 2339 1831 2355
rect 1865 2345 1899 2359
rect 1944 2358 3582 2359
rect 1721 2333 1797 2339
rect 1725 2331 1797 2333
rect 1944 2336 2664 2358
rect 2844 2353 3582 2358
rect 3613 2360 3688 2379
rect 3692 2362 3701 2383
rect 12720 2382 13110 2383
rect 1944 2334 2726 2336
rect 1944 2329 2681 2334
rect 2720 2329 2726 2334
rect 2844 2333 3609 2353
rect 2844 2330 2957 2333
rect 3045 2330 3087 2333
rect 3045 2329 3075 2330
rect 3121 2329 3191 2333
rect 3209 2329 3283 2333
rect 3291 2329 3609 2333
rect 1208 2311 1337 2329
rect 1443 2315 1517 2329
rect 1237 2307 1271 2311
rect 1439 2299 1517 2315
rect 1583 2323 1657 2329
rect 1583 2318 1667 2323
rect 1583 2299 1657 2318
rect 1439 2295 1491 2299
rect 1691 2297 1797 2329
rect 1846 2319 1862 2323
rect 1881 2319 1915 2329
rect 1944 2324 2957 2329
rect 1944 2319 2681 2324
rect 2720 2322 2726 2324
rect 1831 2295 2681 2319
rect 2810 2296 2957 2324
rect 2985 2313 3019 2329
rect 3045 2317 3111 2329
rect 3121 2317 3203 2329
rect 3209 2324 3609 2329
rect 3209 2323 3333 2324
rect 3045 2313 3113 2317
rect 2985 2311 3113 2313
rect 3121 2311 3155 2317
rect 3169 2315 3203 2317
rect 3221 2315 3259 2323
rect 3169 2311 3259 2315
rect 3261 2311 3333 2323
rect 3353 2318 3609 2324
rect 3613 2318 3647 2360
rect 2985 2309 3337 2311
rect 3019 2307 3337 2309
rect 3353 2307 3688 2318
rect 1906 2285 2681 2295
rect 1439 2261 1457 2281
rect 1831 2261 2681 2285
rect 3019 2295 3688 2307
rect 3019 2293 3371 2295
rect 3382 2294 3688 2295
rect 3383 2293 3688 2294
rect 3019 2271 3688 2293
rect 3015 2263 3688 2271
rect 1906 2253 2681 2261
rect 1906 2216 2627 2253
rect 2634 2216 2681 2253
rect 2999 2237 3015 2263
rect 3019 2240 3688 2263
rect 3019 2239 3681 2240
rect 3019 2237 3663 2239
rect 2726 2216 2806 2229
rect 2868 2224 2892 2228
rect 2902 2224 2926 2237
rect 3015 2234 3663 2237
rect 1388 2214 2806 2216
rect 1388 2213 2758 2214
rect 1388 2209 1470 2213
rect 1955 2209 1985 2213
rect 1989 2209 2758 2213
rect 1388 2166 1489 2209
rect 1517 2175 1581 2209
rect 1609 2175 1673 2209
rect 1701 2175 1765 2209
rect 1793 2175 1857 2209
rect 1885 2175 1949 2209
rect 1977 2200 2758 2209
rect 2931 2203 2965 2233
rect 3015 2229 3734 2234
rect 3019 2209 3734 2229
rect 1977 2189 2047 2200
rect 2066 2195 2758 2200
rect 3019 2199 3537 2209
rect 1977 2176 2041 2189
rect 2066 2180 2806 2195
rect 2066 2176 2758 2180
rect 1977 2175 2758 2176
rect 1142 2161 1489 2166
rect 1547 2161 1581 2175
rect 1639 2161 1673 2175
rect 1731 2161 1765 2175
rect 1823 2161 1857 2175
rect 1915 2174 1949 2175
rect 2007 2174 2758 2175
rect 1900 2168 1951 2174
rect 1900 2161 1962 2168
rect 1985 2161 2758 2174
rect 2927 2165 2961 2195
rect 3007 2185 3537 2199
rect 3541 2195 3734 2209
rect 3560 2186 3720 2195
rect 3560 2185 3731 2186
rect 3007 2169 3731 2185
rect 1142 2144 1470 2161
rect 1388 2138 1470 2144
rect 1951 2157 1964 2161
rect 2014 2158 2047 2161
rect 2066 2158 2758 2161
rect 1951 2151 1978 2157
rect 1951 2140 1985 2151
rect 2014 2150 2758 2158
rect 2981 2161 3731 2169
rect 2028 2144 2758 2150
rect 2942 2153 2972 2157
rect 1142 2116 1470 2138
rect 1934 2138 1996 2140
rect 2028 2138 2635 2144
rect 1934 2127 2635 2138
rect 1900 2123 1930 2127
rect 1934 2123 1985 2127
rect 1228 2088 1470 2116
rect 1913 2117 1990 2123
rect 2028 2119 2635 2127
rect 2638 2127 2664 2144
rect 2638 2120 2760 2127
rect 1913 2105 2019 2117
rect 1913 2097 1990 2105
rect 1388 2060 1470 2088
rect 1896 2089 1990 2097
rect 1896 2077 1947 2089
rect 1200 2052 1678 2060
rect 1913 2058 1947 2077
rect 1951 2079 1985 2089
rect 2028 2079 2615 2119
rect 2780 2094 2812 2110
rect 2814 2094 2846 2144
rect 2942 2131 2977 2153
rect 2943 2127 2977 2131
rect 2981 2135 3762 2161
rect 2981 2129 3765 2135
rect 1951 2070 2615 2079
rect 2626 2084 2846 2094
rect 2942 2093 2972 2103
rect 2626 2070 2838 2084
rect 1951 2058 2838 2070
rect 1902 2056 2838 2058
rect 1902 2052 2615 2056
rect 1388 2032 1470 2052
rect 1913 2047 1947 2052
rect 1914 2037 1947 2047
rect 1951 2045 2615 2052
rect 2839 2047 2931 2083
rect 2943 2059 2972 2093
rect 2981 2070 3495 2129
rect 3505 2127 3765 2129
rect 3498 2097 3765 2127
rect 3505 2091 3765 2097
rect 3503 2070 3510 2091
rect 3511 2072 3765 2091
rect 3511 2071 3696 2072
rect 3522 2070 3696 2071
rect 2981 2055 3696 2070
rect 2969 2047 3696 2055
rect 1228 2024 1678 2032
rect 1370 2001 1678 2024
rect 1370 1996 1688 2001
rect 1527 1993 1535 1996
rect 1472 1937 1473 1982
rect 1475 1967 1548 1993
rect 1625 1991 1688 1996
rect 1625 1967 1659 1991
rect 1663 1967 1688 1991
rect 1697 1967 1722 2035
rect 1913 2030 1947 2037
rect 2028 2040 2615 2045
rect 2028 2038 2626 2040
rect 2028 2032 2838 2038
rect 1976 2030 2838 2032
rect 2942 2030 3696 2047
rect 1902 2000 2838 2030
rect 2931 2029 3696 2030
rect 2893 2007 3696 2029
rect 3718 2033 3765 2072
rect 3718 2007 3752 2033
rect 1902 1996 2620 2000
rect 1527 1963 1535 1967
rect 1575 1963 1594 1967
rect 1475 1937 1514 1959
rect 1569 1952 1594 1963
rect 1575 1937 1594 1952
rect 1609 1937 1628 1967
rect 1044 1746 1239 1894
rect 1322 1892 1338 1936
rect 1350 1892 1366 1936
rect 1457 1933 1641 1937
rect 1709 1933 1722 1967
rect 1914 1935 1947 1996
rect 1948 1973 1981 1996
rect 1990 1975 2620 1996
rect 2631 1991 2635 2000
rect 2696 1998 2712 1999
rect 2666 1983 2712 1998
rect 1990 1974 2577 1975
rect 1948 1969 1982 1973
rect 1990 1969 2620 1974
rect 1948 1949 2620 1969
rect 2662 1965 2712 1983
rect 2893 1985 3752 2007
rect 2893 1983 3457 1985
rect 2780 1970 2850 1974
rect 2726 1964 2746 1966
rect 1990 1941 2620 1949
rect 2666 1945 2746 1964
rect 2780 1949 2881 1970
rect 2641 1941 2746 1945
rect 1990 1935 2746 1941
rect 1457 1930 1485 1933
rect 1513 1930 1641 1933
rect 1411 1907 1641 1930
rect 1914 1931 2746 1935
rect 2780 1936 2816 1940
rect 1914 1926 2675 1931
rect 1914 1915 2619 1926
rect 1968 1913 2619 1915
rect 1939 1912 2619 1913
rect 1767 1910 1852 1911
rect 1396 1898 1641 1907
rect 1396 1883 1539 1898
rect 1396 1873 1413 1883
rect 1400 1857 1407 1873
rect 1434 1863 1539 1883
rect 1544 1873 1641 1898
rect 1757 1894 1852 1910
rect 1928 1907 2619 1912
rect 2632 1911 2675 1926
rect 2780 1915 2881 1936
rect 2893 1922 2903 1983
rect 2930 1949 3457 1983
rect 2923 1936 3457 1949
rect 3467 1973 3752 1985
rect 3467 1947 3696 1973
rect 2930 1933 3457 1936
rect 2939 1922 3457 1933
rect 2675 1907 2695 1911
rect 1357 1765 1419 1857
rect 1431 1855 1543 1863
rect 1544 1855 1594 1873
rect 1431 1849 1594 1855
rect 1431 1840 1496 1849
rect 1431 1837 1485 1840
rect 1515 1837 1594 1849
rect 1441 1823 1502 1837
rect 1441 1807 1453 1823
rect 1472 1817 1502 1823
rect 1525 1833 1595 1837
rect 1444 1791 1453 1795
rect 1472 1791 1513 1817
rect 1525 1799 1597 1833
rect 1515 1791 1597 1799
rect 1599 1791 1628 1873
rect 1675 1833 1686 1836
rect 1709 1833 1720 1870
rect 1651 1801 1739 1833
rect 1634 1791 1739 1801
rect 1770 1791 1801 1873
rect 1844 1843 1852 1894
rect 1915 1883 2701 1907
rect 1915 1873 1971 1883
rect 1973 1877 2701 1883
rect 1973 1873 2622 1877
rect 1863 1843 1869 1873
rect 1915 1870 1973 1873
rect 1990 1870 2581 1873
rect 1915 1869 2581 1870
rect 1874 1853 1902 1869
rect 1915 1855 1949 1869
rect 1939 1853 1944 1855
rect 1916 1843 1944 1853
rect 1952 1843 2559 1869
rect 1829 1839 1872 1843
rect 1804 1828 1872 1839
rect 1879 1841 2559 1843
rect 2561 1865 2562 1869
rect 2561 1841 2588 1865
rect 1879 1839 2588 1841
rect 2595 1843 2622 1873
rect 2631 1873 2701 1877
rect 2750 1873 2780 1911
rect 2788 1873 2845 1897
rect 2847 1873 2885 1907
rect 2893 1886 3457 1922
rect 3484 1930 3696 1947
rect 3484 1928 3682 1930
rect 3484 1907 3658 1928
rect 3484 1904 3689 1907
rect 3484 1886 3644 1904
rect 2893 1873 3644 1886
rect 3684 1873 3689 1904
rect 2631 1869 2667 1873
rect 2675 1869 2699 1873
rect 2704 1869 2733 1873
rect 2631 1855 2665 1869
rect 2641 1843 2665 1855
rect 2674 1843 2733 1869
rect 2738 1869 2780 1873
rect 2738 1856 2767 1869
rect 2782 1863 2812 1869
rect 2738 1843 2770 1856
rect 2788 1843 2811 1863
rect 2847 1850 2881 1873
rect 2847 1843 2890 1850
rect 2893 1843 3689 1873
rect 2595 1839 2733 1843
rect 1879 1837 2571 1839
rect 1804 1791 1835 1828
rect 1844 1791 1872 1828
rect 1897 1828 2571 1837
rect 1897 1807 1903 1828
rect 1916 1821 2571 1828
rect 2620 1828 2674 1839
rect 2620 1823 2667 1828
rect 2675 1827 2733 1839
rect 2735 1841 3689 1843
rect 2735 1831 2879 1841
rect 2881 1831 3689 1841
rect 2738 1828 2879 1831
rect 2738 1827 2848 1828
rect 1916 1807 2590 1821
rect 2620 1811 2643 1823
rect 2675 1821 2848 1827
rect 2853 1827 2879 1828
rect 2853 1825 2866 1827
rect 2675 1813 2856 1821
rect 2620 1807 2659 1811
rect 1897 1799 2590 1807
rect 1897 1797 2609 1799
rect 2613 1797 2659 1807
rect 2675 1797 2782 1813
rect 2788 1807 2811 1813
rect 2822 1807 2856 1813
rect 2858 1807 2866 1825
rect 2892 1808 3689 1831
rect 3718 1848 3752 1973
rect 3718 1808 3743 1848
rect 2847 1805 2873 1807
rect 2856 1797 2873 1805
rect 2892 1797 3743 1808
rect 1897 1791 2670 1797
rect 2675 1796 2770 1797
rect 2675 1791 2739 1796
rect 2858 1792 2873 1797
rect 2905 1792 3743 1797
rect 2858 1791 3743 1792
rect 1427 1786 3743 1791
rect 1427 1784 3644 1786
rect 3655 1784 3743 1786
rect 1427 1765 3774 1784
rect 1357 1760 3774 1765
rect 1357 1755 3617 1760
rect 1055 1745 1239 1746
rect 1166 1736 1239 1745
rect 1190 1701 1239 1736
rect 1278 1695 1307 1739
rect 1312 1729 1368 1739
rect 1385 1736 3617 1755
rect 1377 1729 3617 1736
rect 3618 1752 3774 1760
rect 3618 1729 3788 1752
rect 1377 1709 3788 1729
rect 1341 1695 1368 1705
rect 1398 1698 3788 1709
rect 1296 1685 1307 1695
rect 1330 1693 1341 1695
rect 1427 1693 3788 1698
rect 1330 1685 3788 1693
rect 1274 1684 3788 1685
rect 1246 1658 1258 1678
rect 1246 1640 1262 1658
rect 1274 1655 3774 1684
rect 1274 1643 1391 1655
rect 1421 1653 1766 1655
rect 1772 1653 1810 1655
rect 1421 1643 1810 1653
rect 1914 1652 2534 1655
rect 1914 1651 2563 1652
rect 2636 1651 2666 1655
rect 2670 1651 2704 1655
rect 2733 1651 2750 1655
rect 2767 1651 2812 1655
rect 2854 1654 3774 1655
rect 2854 1653 3776 1654
rect 2858 1651 3381 1653
rect 3408 1651 3776 1653
rect 1274 1642 1810 1643
rect 1274 1640 1798 1642
rect 1236 1630 1798 1640
rect 1236 1617 1813 1630
rect 1816 1628 1889 1651
rect 1823 1625 1889 1628
rect 1914 1632 2625 1651
rect 1914 1625 2628 1632
rect 1823 1622 2628 1625
rect 2651 1630 2717 1651
rect 2743 1634 2812 1651
rect 2818 1645 3381 1651
rect 3387 1650 3776 1651
rect 3387 1645 3788 1650
rect 2818 1643 3788 1645
rect 2818 1634 3381 1643
rect 2651 1623 2719 1630
rect 2636 1622 2719 1623
rect 1823 1617 2742 1622
rect 2743 1617 3381 1634
rect 3387 1617 3788 1643
rect 1239 1615 1813 1617
rect 1834 1615 2742 1617
rect 1239 1606 1797 1615
rect 1236 1528 1719 1606
rect 1742 1585 1797 1606
rect 1834 1597 2551 1615
rect 2556 1601 2582 1615
rect 2584 1609 2742 1615
rect 2744 1615 3381 1617
rect 2744 1609 2812 1615
rect 2584 1603 2812 1609
rect 2828 1603 2854 1615
rect 2584 1601 2816 1603
rect 2555 1597 2816 1601
rect 1834 1595 2816 1597
rect 1834 1593 1894 1595
rect 1914 1593 2816 1595
rect 1834 1585 2816 1593
rect 1742 1569 1776 1585
rect 1787 1569 1800 1585
rect 1827 1581 2742 1585
rect 1827 1577 1873 1581
rect 1725 1555 1793 1569
rect 1827 1567 1834 1577
rect 1839 1567 1873 1577
rect 1893 1574 2742 1581
rect 2744 1574 2821 1585
rect 1893 1567 2821 1574
rect 1827 1555 1868 1567
rect 1893 1559 2582 1567
rect 1895 1555 2582 1559
rect 2584 1555 2821 1567
rect 2867 1577 3381 1615
rect 3408 1592 3788 1617
rect 3408 1584 3776 1592
rect 3904 1590 3946 1604
rect 3408 1578 3613 1584
rect 3617 1578 3651 1584
rect 3408 1577 3662 1578
rect 2867 1561 3662 1577
rect 3904 1562 3946 1576
rect 2867 1555 3381 1561
rect 1725 1551 1796 1555
rect 1826 1553 3381 1555
rect 3408 1558 3662 1561
rect 3408 1553 3610 1558
rect 1826 1551 2877 1553
rect 1734 1540 1796 1551
rect 1742 1528 1796 1540
rect 1236 1509 1704 1528
rect 1734 1509 1796 1528
rect 1236 1503 1796 1509
rect 1821 1523 2816 1551
rect 1821 1513 1827 1523
rect 1840 1519 2816 1523
rect 2820 1545 2877 1551
rect 2982 1549 2986 1551
rect 3020 1549 3110 1553
rect 3112 1549 3144 1553
rect 3148 1551 3174 1553
rect 3182 1551 3201 1553
rect 3204 1551 3279 1553
rect 3148 1549 3279 1551
rect 3283 1549 3381 1553
rect 3382 1549 3610 1553
rect 2893 1547 2927 1549
rect 2982 1547 3610 1549
rect 2893 1545 2903 1547
rect 2954 1545 3610 1547
rect 2820 1531 2933 1545
rect 2954 1538 3020 1545
rect 1840 1515 2774 1519
rect 1840 1513 1894 1515
rect 1821 1503 1894 1513
rect 1914 1508 2774 1515
rect 1921 1506 2035 1508
rect 2036 1506 2774 1508
rect 1921 1503 2774 1506
rect 2782 1517 2790 1519
rect 2820 1517 2957 1531
rect 2982 1527 3020 1538
rect 2782 1503 2797 1517
rect 2816 1509 2957 1517
rect 2820 1503 2957 1509
rect 2983 1503 2986 1515
rect 3017 1503 3020 1515
rect 3023 1503 3053 1545
rect 3061 1529 3610 1545
rect 3613 1541 3651 1548
rect 3061 1520 3613 1529
rect 3061 1505 3712 1520
rect 3718 1505 3740 1548
rect 3994 1536 4070 1544
rect 3880 1505 3904 1530
rect 3908 1505 3932 1530
rect 4146 1520 4170 1528
rect 3966 1508 4042 1516
rect 3061 1503 3666 1505
rect 1236 1498 3666 1503
rect 1236 1496 3578 1498
rect 3579 1496 3666 1498
rect 1198 1472 3666 1496
rect 1198 1461 3541 1472
rect 1198 1441 1300 1461
rect 1301 1441 3541 1461
rect 3542 1441 3666 1472
rect 1198 1417 3666 1441
rect 1198 1407 1300 1417
rect 1320 1408 3666 1417
rect 1198 1388 1305 1407
rect 1330 1397 1339 1408
rect 1351 1405 3666 1408
rect 1200 1364 1224 1388
rect 1254 1386 1305 1388
rect 1258 1383 1305 1386
rect 1345 1393 3666 1405
rect 1286 1374 1339 1383
rect 1296 1363 1339 1374
rect 1345 1376 3540 1393
rect 3542 1385 3666 1393
rect 1345 1359 1350 1376
rect 1351 1367 3540 1376
rect 1358 1365 1666 1367
rect 1696 1365 1758 1367
rect 1358 1363 1758 1365
rect 1783 1363 1789 1367
rect 1802 1363 1856 1367
rect 1883 1363 1997 1367
rect 1998 1363 2021 1367
rect 2035 1363 2107 1367
rect 1358 1359 1997 1363
rect 2023 1359 2107 1363
rect 2115 1364 2458 1367
rect 2461 1364 2560 1367
rect 2115 1359 2560 1364
rect 2595 1365 2668 1367
rect 2595 1363 2628 1365
rect 2706 1363 2736 1367
rect 2575 1359 2641 1363
rect 2667 1359 2736 1363
rect 2744 1359 2919 1367
rect 2928 1366 3540 1367
rect 3541 1366 3666 1385
rect 2928 1362 3666 1366
rect 3682 1496 3932 1505
rect 2928 1361 3647 1362
rect 2928 1360 3629 1361
rect 3682 1360 3712 1496
rect 2928 1359 3712 1360
rect 1313 1354 3712 1359
rect 1244 1297 1261 1331
rect 1263 1328 3712 1354
rect 1263 1297 3628 1328
rect 1254 1273 3628 1297
rect 3682 1304 3712 1328
rect 3718 1304 3740 1496
rect 3880 1412 3904 1496
rect 3908 1412 3932 1496
rect 3956 1392 4032 1400
rect 8902 1378 9106 1380
rect 3928 1364 4004 1372
rect 3682 1296 3700 1304
rect 3718 1278 3720 1304
rect 1282 1270 3628 1273
rect 1186 1264 3628 1270
rect 3842 1268 3866 1302
rect 3870 1268 3894 1302
rect 1220 1242 1267 1263
rect 1270 1258 3628 1264
rect 1292 1253 1301 1258
rect 1307 1249 3628 1258
rect 1307 1242 3502 1249
rect 1186 1236 3502 1242
rect 1242 1230 3502 1236
rect 1258 1219 1301 1230
rect 1307 1215 1312 1230
rect 1313 1223 3502 1230
rect 1320 1221 1628 1223
rect 1658 1221 1720 1223
rect 1320 1219 1720 1221
rect 1745 1219 1751 1223
rect 1764 1219 1818 1223
rect 1320 1215 1743 1219
rect 1764 1215 1835 1219
rect 1845 1215 1959 1223
rect 1960 1219 1983 1223
rect 1997 1219 2698 1223
rect 1967 1215 2698 1219
rect 2706 1215 2881 1223
rect 2907 1219 2910 1223
rect 2928 1215 2984 1223
rect 2985 1222 3502 1223
rect 3504 1222 3628 1249
rect 3918 1248 3994 1256
rect 2985 1218 3628 1222
rect 3890 1220 3966 1228
rect 2985 1217 3609 1218
rect 2985 1216 3591 1217
rect 2985 1215 3644 1216
rect 1275 1211 3644 1215
rect 1231 1210 3644 1211
rect 1225 1184 3644 1210
rect 1225 1163 3590 1184
rect 1232 1147 3590 1163
rect 1233 1145 3590 1147
rect 1244 1132 3590 1145
rect 1210 1120 1238 1129
rect 1244 1128 3628 1132
rect 3828 1128 3832 1152
rect 8196 1150 8224 1152
rect 1244 1120 3590 1128
rect 3804 1124 3828 1128
rect 3832 1124 3856 1128
rect 1210 1114 3590 1120
rect 1210 1095 1250 1114
rect 1254 1109 3590 1114
rect 1262 1104 3590 1109
rect 1262 1100 3628 1104
rect 3828 1100 3832 1124
rect 3880 1104 3956 1112
rect 1262 1095 3464 1100
rect 1210 1091 3464 1095
rect 1216 1088 3464 1091
rect 3466 1088 3590 1100
rect 1216 1086 3590 1088
rect 1220 1079 3590 1086
rect 1220 1075 1429 1079
rect 1262 1071 1429 1075
rect 1539 1071 1722 1079
rect 1728 1078 1780 1079
rect 1783 1078 1890 1079
rect 1728 1075 1890 1078
rect 1920 1075 1977 1079
rect 1728 1071 1794 1075
rect 1807 1071 1981 1075
rect 1997 1071 2103 1079
rect 2115 1075 2137 1079
rect 2139 1075 2418 1079
rect 2115 1071 2418 1075
rect 2423 1071 2442 1079
rect 2458 1075 2475 1079
rect 2492 1077 3590 1079
rect 2492 1075 2630 1077
rect 2475 1071 2630 1075
rect 2660 1074 3590 1077
rect 3852 1076 3928 1084
rect 2660 1073 3571 1074
rect 2660 1072 3458 1073
rect 2660 1071 3444 1072
rect 1237 1066 3444 1071
rect 1183 1063 3444 1066
rect 1220 990 1232 1035
rect 1237 1031 3444 1063
rect 3518 1040 3606 1072
rect 4006 1068 4032 1072
rect 4034 1040 4060 1072
rect 1237 1029 2766 1031
rect 1237 1007 2796 1029
rect 2833 1028 3044 1031
rect 3074 1028 3220 1031
rect 2833 1010 3220 1028
rect 2833 1007 2953 1010
rect 1237 990 2766 1007
rect 1208 970 2766 990
rect 2878 985 2879 1007
rect 1220 969 1232 970
rect 1157 965 1232 969
rect 1237 965 2766 970
rect 1157 961 2766 965
rect 2895 983 2953 1007
rect 2962 1004 3128 1010
rect 3165 1007 3220 1010
rect 3170 1004 3220 1007
rect 2962 1003 3220 1004
rect 2895 961 2947 983
rect 2962 961 3044 1003
rect 3074 990 3220 1003
rect 3244 990 3248 1031
rect 3250 1001 3296 1031
rect 3250 990 3304 1001
rect 3334 990 3396 1001
rect 3074 982 3396 990
rect 3074 961 3136 982
rect 3146 980 3396 982
rect 3146 962 3220 980
rect 3244 976 3248 980
rect 3250 976 3320 980
rect 3250 962 3304 976
rect 3334 962 3396 980
rect 3146 961 3402 962
rect 1157 955 2789 961
rect 882 902 909 911
rect 910 902 937 939
rect 1157 931 1232 955
rect 1236 954 2789 955
rect 1236 953 2747 954
rect 1236 952 2634 953
rect 1236 943 2620 952
rect 2645 943 2713 953
rect 1236 942 2713 943
rect 1237 939 2713 942
rect 1237 935 2620 939
rect 1239 931 1528 935
rect 1157 927 1528 931
rect 1541 927 1575 931
rect 1578 927 1897 935
rect 1927 931 2065 935
rect 1921 927 2065 931
rect 2075 927 2085 935
rect 2097 931 2346 935
rect 2093 927 2346 931
rect 2358 927 2385 935
rect 2437 931 2620 935
rect 2442 927 2620 931
rect 1157 911 2620 927
rect 2645 923 2713 939
rect 2721 935 2740 953
rect 2759 935 2789 954
rect 2947 949 2987 961
rect 2947 947 2977 949
rect 3006 947 3019 961
rect 3044 947 3074 961
rect 3098 947 3116 961
rect 3136 952 3402 961
rect 3136 947 3166 952
rect 3176 947 3208 952
rect 3220 947 3250 952
rect 3266 947 3292 952
rect 3304 947 3350 952
rect 2947 935 2992 947
rect 1277 901 1304 911
rect 1317 901 1349 911
rect 1541 901 1575 911
rect 1579 901 1613 905
rect 1616 901 1651 911
rect 1681 901 1793 911
rect 1225 897 1277 901
rect 1307 897 1399 901
rect 1513 899 1651 901
rect 1225 887 1361 897
rect 1225 874 1303 887
rect 1307 886 1361 887
rect 1225 866 1308 874
rect 1225 863 1303 866
rect 1317 863 1361 886
rect 1225 851 1367 863
rect 1225 846 1327 851
rect 1216 838 1327 846
rect 1225 825 1327 838
rect 1207 821 1327 825
rect 1164 817 1327 821
rect 1164 803 1329 817
rect 1277 791 1293 803
rect 1301 791 1329 803
rect 1301 787 1327 791
rect 1343 787 1367 851
rect 1395 817 1401 889
rect 1433 839 1435 897
rect 1437 817 1443 879
rect 1467 821 1469 897
rect 1513 886 1528 899
rect 1533 897 1651 899
rect 1677 899 1793 901
rect 1795 899 1851 911
rect 1921 901 1943 911
rect 1677 897 1851 899
rect 1855 897 1943 901
rect 2001 901 2035 911
rect 2044 901 2045 911
rect 2093 901 2103 911
rect 2104 901 2177 911
rect 2001 899 2177 901
rect 2001 897 2045 899
rect 1533 889 1643 897
rect 1549 887 1643 889
rect 1475 821 1481 841
rect 1511 832 1547 879
rect 1561 865 1643 887
rect 1647 865 1675 897
rect 1677 889 1696 897
rect 1795 889 1829 897
rect 1855 891 1952 897
rect 1837 889 1952 891
rect 1677 886 1952 889
rect 2029 886 2045 897
rect 1677 874 1883 886
rect 1677 865 1787 874
rect 1795 871 1883 874
rect 1897 871 1927 886
rect 1795 866 1929 871
rect 1561 863 1647 865
rect 1677 863 1795 865
rect 1561 855 1643 863
rect 1561 839 1615 855
rect 1681 843 1711 863
rect 1561 835 1591 839
rect 1657 835 1711 843
rect 1715 857 1787 863
rect 1801 857 1807 866
rect 1811 857 1883 866
rect 1715 843 1855 857
rect 1897 843 1927 866
rect 1715 838 1927 843
rect 1715 835 1855 838
rect 1897 835 1927 838
rect 1937 835 1952 886
rect 2044 849 2045 886
rect 2054 865 2177 899
rect 2185 908 2261 911
rect 2185 897 2266 908
rect 2277 897 2304 911
rect 2075 849 2177 865
rect 2085 835 2115 849
rect 1561 832 2130 835
rect 1377 787 1401 817
rect 1467 791 1507 821
rect 1511 817 2130 832
rect 2167 821 2172 849
rect 2201 825 2206 897
rect 2207 889 2266 897
rect 2346 889 2348 911
rect 2390 899 2424 911
rect 2458 901 2471 911
rect 2481 909 2560 911
rect 2481 901 2611 909
rect 2431 899 2481 901
rect 2390 897 2481 899
rect 2505 897 2611 901
rect 2645 897 2679 923
rect 2737 897 2751 931
rect 2954 920 2969 935
rect 2977 932 2992 935
rect 3036 935 3089 947
rect 3036 932 3044 935
rect 3074 932 3089 935
rect 3128 935 3206 947
rect 3128 932 3136 935
rect 3138 933 3206 935
rect 3142 932 3206 933
rect 3212 935 3265 947
rect 3212 932 3220 935
rect 3250 932 3265 935
rect 3296 935 3350 947
rect 3296 932 3304 935
rect 3142 931 3172 932
rect 3176 931 3206 932
rect 3320 931 3350 935
rect 3354 931 3384 952
rect 2915 897 3030 913
rect 2207 849 2276 889
rect 2331 877 2390 889
rect 2415 877 2492 897
rect 3480 896 3568 928
rect 3766 896 3790 1014
rect 3794 924 3818 1014
rect 2331 874 2472 877
rect 2346 865 2472 874
rect 2346 849 2385 865
rect 2390 863 2472 865
rect 2415 849 2472 863
rect 2539 863 2577 875
rect 2949 863 2996 879
rect 2207 827 2212 849
rect 2274 827 2276 849
rect 2221 825 2255 827
rect 2315 821 2424 849
rect 2442 827 2472 849
rect 2505 827 2526 855
rect 1573 791 1613 817
rect 1616 791 1633 817
rect 1657 813 1688 817
rect 1715 813 1821 817
rect 1657 791 1687 813
rect 1711 797 1821 813
rect 1855 803 1889 817
rect 1937 797 1952 817
rect 1711 791 1787 797
rect 2085 793 2115 817
rect 2159 793 2172 821
rect 2442 817 2457 827
rect 1715 789 1787 791
rect 2059 791 2125 793
rect 2177 791 2182 817
rect 2304 791 2306 817
rect 2388 815 2415 817
rect 2059 787 2091 791
rect 2093 787 2125 791
rect 2314 787 2348 815
rect 2382 787 2424 815
rect 2481 791 2526 827
rect 2505 787 2526 791
rect 2539 787 2560 863
rect 2564 817 2630 852
rect 2660 845 2751 852
rect 2660 817 2764 845
rect 8902 834 8907 868
rect 8902 833 8941 834
rect 2618 792 2710 798
rect 2619 791 2671 792
rect 2619 787 2630 791
rect 2660 787 2671 791
rect 1198 769 1327 787
rect 1433 773 1507 787
rect 1227 765 1261 769
rect 1429 757 1507 773
rect 1573 781 1647 787
rect 1573 776 1657 781
rect 1573 757 1647 776
rect 1429 753 1481 757
rect 1681 755 1787 787
rect 1836 777 1852 781
rect 1871 777 1905 787
rect 1821 753 1937 777
rect 1958 776 1979 781
rect 2033 776 2085 781
rect 2091 759 2093 787
rect 2159 759 2206 787
rect 1429 726 1447 739
rect 1821 726 1937 743
rect 1198 724 2610 726
rect 1198 722 2728 724
rect 1429 719 1447 722
rect 1821 719 1937 722
rect 1170 696 2582 698
rect 1170 694 2728 696
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use cp_schem  cp_schem_0
timestamp 1708425511
transform 1 0 5618 0 1 2600
box 1298 4024 6324 5767
use cp_schem  cp_schem_1
timestamp 1708425511
transform 1 0 5656 0 1 2600
box 1298 4024 6324 5767
use cp_schem  cp_schem_2
timestamp 1708425511
transform 1 0 5694 0 1 2600
box 1298 4024 6324 5767
use cp_schem  cp_schem_3
timestamp 1708425511
transform 1 0 5732 0 1 2600
box 1298 4024 6324 5767
use cp_schem  cp_schem_4
timestamp 1708425511
transform 1 0 5770 0 1 2600
box 1298 4024 6324 5767
use cp_schem  cp_schem_5
timestamp 1708425511
transform 1 0 5846 0 1 2600
box 1298 4024 6324 5767
use cp_schem  cp_schem_6
timestamp 1708425511
transform 1 0 -1298 0 1 -6024
box 1298 4024 6324 5767
use inverter  inverter_0
timestamp 1708425308
transform 1 0 12222 0 1 1800
box -280 -1200 1040 1362
use inverter  inverter_1
timestamp 1708425308
transform 1 0 12260 0 1 1800
box -280 -1200 1040 1362
use inverter  inverter_2
timestamp 1708425308
transform 1 0 12298 0 1 1800
box -280 -1200 1040 1362
use inverter  inverter_3
timestamp 1708425308
transform 1 0 12336 0 1 1800
box -280 -1200 1040 1362
use inverter  inverter_4
timestamp 1708425308
transform 1 0 12374 0 1 1800
box -280 -1200 1040 1362
use inverter  inverter_5
timestamp 1708425308
transform 1 0 12450 0 1 1800
box -280 -1200 1040 1362
use inverter  inverter_6
timestamp 1708425308
transform 1 0 5306 0 1 -800
box -280 -1200 1040 1362
use pfd  pfd_0
timestamp 1708426743
transform 1 0 38 0 1 2600
box 786 -1880 3956 334
use pfd  pfd_1
timestamp 1708426743
transform 1 0 76 0 1 2744
box 786 -1880 3956 334
use pfd  pfd_2
timestamp 1708426743
transform 1 0 114 0 1 2888
box 786 -1880 3956 334
use pfd  pfd_3
timestamp 1708426743
transform 1 0 152 0 1 3032
box 786 -1880 3956 334
use pfd  pfd_4
timestamp 1708426743
transform 1 0 190 0 1 3176
box 786 -1880 3956 334
use pfd  pfd_5
timestamp 1708426743
transform 1 0 266 0 1 3464
box 786 -1880 3956 334
use pfd  x1
timestamp 1708426743
transform 1 0 -786 0 1 2480
box 786 -1880 3956 334
use cp_schem  x2
timestamp 1708425511
transform 1 0 1872 0 1 -3424
box 1298 4024 6324 5767
use inverter  x3
timestamp 1708425308
transform 1 0 8476 0 1 216
box -280 -1200 1040 1362
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 cp_bias
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 cp_out
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 B
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
