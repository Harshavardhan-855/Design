magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< error_p >>
rect -560 154 -502 160
rect -442 154 -384 160
rect -324 154 -266 160
rect -206 154 -148 160
rect -88 154 -30 160
rect 30 154 88 160
rect 148 154 206 160
rect 266 154 324 160
rect 384 154 442 160
rect 502 154 560 160
rect -560 120 -548 154
rect -442 120 -430 154
rect -324 120 -312 154
rect -206 120 -194 154
rect -88 120 -76 154
rect 30 120 42 154
rect 148 120 160 154
rect 266 120 278 154
rect 384 120 396 154
rect 502 120 514 154
rect -560 114 -502 120
rect -442 114 -384 120
rect -324 114 -266 120
rect -206 114 -148 120
rect -88 114 -30 120
rect 30 114 88 120
rect 148 114 206 120
rect 266 114 324 120
rect 384 114 442 120
rect 502 114 560 120
rect -560 -120 -502 -114
rect -442 -120 -384 -114
rect -324 -120 -266 -114
rect -206 -120 -148 -114
rect -88 -120 -30 -114
rect 30 -120 88 -114
rect 148 -120 206 -114
rect 266 -120 324 -114
rect 384 -120 442 -114
rect 502 -120 560 -114
rect -560 -154 -548 -120
rect -442 -154 -430 -120
rect -324 -154 -312 -120
rect -206 -154 -194 -120
rect -88 -154 -76 -120
rect 30 -154 42 -120
rect 148 -154 160 -120
rect 266 -154 278 -120
rect 384 -154 396 -120
rect 502 -154 514 -120
rect -560 -160 -502 -154
rect -442 -160 -384 -154
rect -324 -160 -266 -154
rect -206 -160 -148 -154
rect -88 -160 -30 -154
rect 30 -160 88 -154
rect 148 -160 206 -154
rect 266 -160 324 -154
rect 384 -160 442 -154
rect 502 -160 560 -154
<< pwell >>
rect -757 -292 757 292
<< nmos >>
rect -561 -82 -501 82
rect -443 -82 -383 82
rect -325 -82 -265 82
rect -207 -82 -147 82
rect -89 -82 -29 82
rect 29 -82 89 82
rect 147 -82 207 82
rect 265 -82 325 82
rect 383 -82 443 82
rect 501 -82 561 82
<< ndiff >>
rect -619 70 -561 82
rect -619 -70 -607 70
rect -573 -70 -561 70
rect -619 -82 -561 -70
rect -501 70 -443 82
rect -501 -70 -489 70
rect -455 -70 -443 70
rect -501 -82 -443 -70
rect -383 70 -325 82
rect -383 -70 -371 70
rect -337 -70 -325 70
rect -383 -82 -325 -70
rect -265 70 -207 82
rect -265 -70 -253 70
rect -219 -70 -207 70
rect -265 -82 -207 -70
rect -147 70 -89 82
rect -147 -70 -135 70
rect -101 -70 -89 70
rect -147 -82 -89 -70
rect -29 70 29 82
rect -29 -70 -17 70
rect 17 -70 29 70
rect -29 -82 29 -70
rect 89 70 147 82
rect 89 -70 101 70
rect 135 -70 147 70
rect 89 -82 147 -70
rect 207 70 265 82
rect 207 -70 219 70
rect 253 -70 265 70
rect 207 -82 265 -70
rect 325 70 383 82
rect 325 -70 337 70
rect 371 -70 383 70
rect 325 -82 383 -70
rect 443 70 501 82
rect 443 -70 455 70
rect 489 -70 501 70
rect 443 -82 501 -70
rect 561 70 619 82
rect 561 -70 573 70
rect 607 -70 619 70
rect 561 -82 619 -70
<< ndiffc >>
rect -607 -70 -573 70
rect -489 -70 -455 70
rect -371 -70 -337 70
rect -253 -70 -219 70
rect -135 -70 -101 70
rect -17 -70 17 70
rect 101 -70 135 70
rect 219 -70 253 70
rect 337 -70 371 70
rect 455 -70 489 70
rect 573 -70 607 70
<< psubdiff >>
rect -721 222 -625 256
rect 625 222 721 256
rect -721 160 -687 222
rect 687 160 721 222
rect -721 -222 -687 -160
rect 687 -222 721 -160
rect -721 -256 -625 -222
rect 625 -256 721 -222
<< psubdiffcont >>
rect -625 222 625 256
rect -721 -160 -687 160
rect 687 -160 721 160
rect -625 -256 625 -222
<< poly >>
rect -564 154 -498 170
rect -564 120 -548 154
rect -514 120 -498 154
rect -564 104 -498 120
rect -446 154 -380 170
rect -446 120 -430 154
rect -396 120 -380 154
rect -446 104 -380 120
rect -328 154 -262 170
rect -328 120 -312 154
rect -278 120 -262 154
rect -328 104 -262 120
rect -210 154 -144 170
rect -210 120 -194 154
rect -160 120 -144 154
rect -210 104 -144 120
rect -92 154 -26 170
rect -92 120 -76 154
rect -42 120 -26 154
rect -92 104 -26 120
rect 26 154 92 170
rect 26 120 42 154
rect 76 120 92 154
rect 26 104 92 120
rect 144 154 210 170
rect 144 120 160 154
rect 194 120 210 154
rect 144 104 210 120
rect 262 154 328 170
rect 262 120 278 154
rect 312 120 328 154
rect 262 104 328 120
rect 380 154 446 170
rect 380 120 396 154
rect 430 120 446 154
rect 380 104 446 120
rect 498 154 564 170
rect 498 120 514 154
rect 548 120 564 154
rect 498 104 564 120
rect -561 82 -501 104
rect -443 82 -383 104
rect -325 82 -265 104
rect -207 82 -147 104
rect -89 82 -29 104
rect 29 82 89 104
rect 147 82 207 104
rect 265 82 325 104
rect 383 82 443 104
rect 501 82 561 104
rect -561 -104 -501 -82
rect -443 -104 -383 -82
rect -325 -104 -265 -82
rect -207 -104 -147 -82
rect -89 -104 -29 -82
rect 29 -104 89 -82
rect 147 -104 207 -82
rect 265 -104 325 -82
rect 383 -104 443 -82
rect 501 -104 561 -82
rect -564 -120 -498 -104
rect -564 -154 -548 -120
rect -514 -154 -498 -120
rect -564 -170 -498 -154
rect -446 -120 -380 -104
rect -446 -154 -430 -120
rect -396 -154 -380 -120
rect -446 -170 -380 -154
rect -328 -120 -262 -104
rect -328 -154 -312 -120
rect -278 -154 -262 -120
rect -328 -170 -262 -154
rect -210 -120 -144 -104
rect -210 -154 -194 -120
rect -160 -154 -144 -120
rect -210 -170 -144 -154
rect -92 -120 -26 -104
rect -92 -154 -76 -120
rect -42 -154 -26 -120
rect -92 -170 -26 -154
rect 26 -120 92 -104
rect 26 -154 42 -120
rect 76 -154 92 -120
rect 26 -170 92 -154
rect 144 -120 210 -104
rect 144 -154 160 -120
rect 194 -154 210 -120
rect 144 -170 210 -154
rect 262 -120 328 -104
rect 262 -154 278 -120
rect 312 -154 328 -120
rect 262 -170 328 -154
rect 380 -120 446 -104
rect 380 -154 396 -120
rect 430 -154 446 -120
rect 380 -170 446 -154
rect 498 -120 564 -104
rect 498 -154 514 -120
rect 548 -154 564 -120
rect 498 -170 564 -154
<< polycont >>
rect -548 120 -514 154
rect -430 120 -396 154
rect -312 120 -278 154
rect -194 120 -160 154
rect -76 120 -42 154
rect 42 120 76 154
rect 160 120 194 154
rect 278 120 312 154
rect 396 120 430 154
rect 514 120 548 154
rect -548 -154 -514 -120
rect -430 -154 -396 -120
rect -312 -154 -278 -120
rect -194 -154 -160 -120
rect -76 -154 -42 -120
rect 42 -154 76 -120
rect 160 -154 194 -120
rect 278 -154 312 -120
rect 396 -154 430 -120
rect 514 -154 548 -120
<< locali >>
rect -721 222 -625 256
rect 625 222 721 256
rect -721 160 -687 222
rect 687 160 721 222
rect -564 120 -548 154
rect -514 120 -498 154
rect -446 120 -430 154
rect -396 120 -380 154
rect -328 120 -312 154
rect -278 120 -262 154
rect -210 120 -194 154
rect -160 120 -144 154
rect -92 120 -76 154
rect -42 120 -26 154
rect 26 120 42 154
rect 76 120 92 154
rect 144 120 160 154
rect 194 120 210 154
rect 262 120 278 154
rect 312 120 328 154
rect 380 120 396 154
rect 430 120 446 154
rect 498 120 514 154
rect 548 120 564 154
rect -607 70 -573 86
rect -607 -86 -573 -70
rect -489 70 -455 86
rect -489 -86 -455 -70
rect -371 70 -337 86
rect -371 -86 -337 -70
rect -253 70 -219 86
rect -253 -86 -219 -70
rect -135 70 -101 86
rect -135 -86 -101 -70
rect -17 70 17 86
rect -17 -86 17 -70
rect 101 70 135 86
rect 101 -86 135 -70
rect 219 70 253 86
rect 219 -86 253 -70
rect 337 70 371 86
rect 337 -86 371 -70
rect 455 70 489 86
rect 455 -86 489 -70
rect 573 70 607 86
rect 573 -86 607 -70
rect -564 -154 -548 -120
rect -514 -154 -498 -120
rect -446 -154 -430 -120
rect -396 -154 -380 -120
rect -328 -154 -312 -120
rect -278 -154 -262 -120
rect -210 -154 -194 -120
rect -160 -154 -144 -120
rect -92 -154 -76 -120
rect -42 -154 -26 -120
rect 26 -154 42 -120
rect 76 -154 92 -120
rect 144 -154 160 -120
rect 194 -154 210 -120
rect 262 -154 278 -120
rect 312 -154 328 -120
rect 380 -154 396 -120
rect 430 -154 446 -120
rect 498 -154 514 -120
rect 548 -154 564 -120
rect -721 -222 -687 -160
rect 687 -222 721 -160
rect -721 -256 -625 -222
rect 625 -256 721 -222
<< viali >>
rect -548 120 -514 154
rect -430 120 -396 154
rect -312 120 -278 154
rect -194 120 -160 154
rect -76 120 -42 154
rect 42 120 76 154
rect 160 120 194 154
rect 278 120 312 154
rect 396 120 430 154
rect 514 120 548 154
rect -607 -70 -573 70
rect -489 -70 -455 70
rect -371 -70 -337 70
rect -253 -70 -219 70
rect -135 -70 -101 70
rect -17 -70 17 70
rect 101 -70 135 70
rect 219 -70 253 70
rect 337 -70 371 70
rect 455 -70 489 70
rect 573 -70 607 70
rect -548 -154 -514 -120
rect -430 -154 -396 -120
rect -312 -154 -278 -120
rect -194 -154 -160 -120
rect -76 -154 -42 -120
rect 42 -154 76 -120
rect 160 -154 194 -120
rect 278 -154 312 -120
rect 396 -154 430 -120
rect 514 -154 548 -120
<< metal1 >>
rect -560 154 -502 160
rect -560 120 -548 154
rect -514 120 -502 154
rect -560 114 -502 120
rect -442 154 -384 160
rect -442 120 -430 154
rect -396 120 -384 154
rect -442 114 -384 120
rect -324 154 -266 160
rect -324 120 -312 154
rect -278 120 -266 154
rect -324 114 -266 120
rect -206 154 -148 160
rect -206 120 -194 154
rect -160 120 -148 154
rect -206 114 -148 120
rect -88 154 -30 160
rect -88 120 -76 154
rect -42 120 -30 154
rect -88 114 -30 120
rect 30 154 88 160
rect 30 120 42 154
rect 76 120 88 154
rect 30 114 88 120
rect 148 154 206 160
rect 148 120 160 154
rect 194 120 206 154
rect 148 114 206 120
rect 266 154 324 160
rect 266 120 278 154
rect 312 120 324 154
rect 266 114 324 120
rect 384 154 442 160
rect 384 120 396 154
rect 430 120 442 154
rect 384 114 442 120
rect 502 154 560 160
rect 502 120 514 154
rect 548 120 560 154
rect 502 114 560 120
rect -613 70 -567 82
rect -613 -70 -607 70
rect -573 -70 -567 70
rect -613 -82 -567 -70
rect -495 70 -449 82
rect -495 -70 -489 70
rect -455 -70 -449 70
rect -495 -82 -449 -70
rect -377 70 -331 82
rect -377 -70 -371 70
rect -337 -70 -331 70
rect -377 -82 -331 -70
rect -259 70 -213 82
rect -259 -70 -253 70
rect -219 -70 -213 70
rect -259 -82 -213 -70
rect -141 70 -95 82
rect -141 -70 -135 70
rect -101 -70 -95 70
rect -141 -82 -95 -70
rect -23 70 23 82
rect -23 -70 -17 70
rect 17 -70 23 70
rect -23 -82 23 -70
rect 95 70 141 82
rect 95 -70 101 70
rect 135 -70 141 70
rect 95 -82 141 -70
rect 213 70 259 82
rect 213 -70 219 70
rect 253 -70 259 70
rect 213 -82 259 -70
rect 331 70 377 82
rect 331 -70 337 70
rect 371 -70 377 70
rect 331 -82 377 -70
rect 449 70 495 82
rect 449 -70 455 70
rect 489 -70 495 70
rect 449 -82 495 -70
rect 567 70 613 82
rect 567 -70 573 70
rect 607 -70 613 70
rect 567 -82 613 -70
rect -560 -120 -502 -114
rect -560 -154 -548 -120
rect -514 -154 -502 -120
rect -560 -160 -502 -154
rect -442 -120 -384 -114
rect -442 -154 -430 -120
rect -396 -154 -384 -120
rect -442 -160 -384 -154
rect -324 -120 -266 -114
rect -324 -154 -312 -120
rect -278 -154 -266 -120
rect -324 -160 -266 -154
rect -206 -120 -148 -114
rect -206 -154 -194 -120
rect -160 -154 -148 -120
rect -206 -160 -148 -154
rect -88 -120 -30 -114
rect -88 -154 -76 -120
rect -42 -154 -30 -120
rect -88 -160 -30 -154
rect 30 -120 88 -114
rect 30 -154 42 -120
rect 76 -154 88 -120
rect 30 -160 88 -154
rect 148 -120 206 -114
rect 148 -154 160 -120
rect 194 -154 206 -120
rect 148 -160 206 -154
rect 266 -120 324 -114
rect 266 -154 278 -120
rect 312 -154 324 -120
rect 266 -160 324 -154
rect 384 -120 442 -114
rect 384 -154 396 -120
rect 430 -154 442 -120
rect 384 -160 442 -154
rect 502 -120 560 -114
rect 502 -154 514 -120
rect 548 -154 560 -120
rect 502 -160 560 -154
<< properties >>
string FIXED_BBOX -704 -239 704 239
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.82 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
