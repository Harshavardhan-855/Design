magic
tech sky130A
magscale 1 2
timestamp 1707817411
<< error_p >>
rect -29 2117 29 2123
rect -29 2083 -17 2117
rect -29 2077 29 2083
rect -29 789 29 795
rect -29 755 -17 789
rect -29 749 29 755
rect -29 681 29 687
rect -29 647 -17 681
rect -29 641 29 647
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect -29 -687 29 -681
rect -29 -755 29 -749
rect -29 -789 -17 -755
rect -29 -795 29 -789
rect -29 -2083 29 -2077
rect -29 -2117 -17 -2083
rect -29 -2123 29 -2117
<< nwell >>
rect -226 -2255 226 2255
<< pmos >>
rect -30 836 30 2036
rect -30 -600 30 600
rect -30 -2036 30 -836
<< pdiff >>
rect -88 2024 -30 2036
rect -88 848 -76 2024
rect -42 848 -30 2024
rect -88 836 -30 848
rect 30 2024 88 2036
rect 30 848 42 2024
rect 76 848 88 2024
rect 30 836 88 848
rect -88 588 -30 600
rect -88 -588 -76 588
rect -42 -588 -30 588
rect -88 -600 -30 -588
rect 30 588 88 600
rect 30 -588 42 588
rect 76 -588 88 588
rect 30 -600 88 -588
rect -88 -848 -30 -836
rect -88 -2024 -76 -848
rect -42 -2024 -30 -848
rect -88 -2036 -30 -2024
rect 30 -848 88 -836
rect 30 -2024 42 -848
rect 76 -2024 88 -848
rect 30 -2036 88 -2024
<< pdiffc >>
rect -76 848 -42 2024
rect 42 848 76 2024
rect -76 -588 -42 588
rect 42 -588 76 588
rect -76 -2024 -42 -848
rect 42 -2024 76 -848
<< nsubdiff >>
rect -190 2185 -94 2219
rect 94 2185 190 2219
rect -190 2123 -156 2185
rect 156 2123 190 2185
rect -190 -2185 -156 -2123
rect 156 -2185 190 -2123
rect -190 -2219 -94 -2185
rect 94 -2219 190 -2185
<< nsubdiffcont >>
rect -94 2185 94 2219
rect -190 -2123 -156 2123
rect 156 -2123 190 2123
rect -94 -2219 94 -2185
<< poly >>
rect -33 2117 33 2133
rect -33 2083 -17 2117
rect 17 2083 33 2117
rect -33 2067 33 2083
rect -30 2036 30 2067
rect -30 805 30 836
rect -33 789 33 805
rect -33 755 -17 789
rect 17 755 33 789
rect -33 739 33 755
rect -33 681 33 697
rect -33 647 -17 681
rect 17 647 33 681
rect -33 631 33 647
rect -30 600 30 631
rect -30 -631 30 -600
rect -33 -647 33 -631
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -697 33 -681
rect -33 -755 33 -739
rect -33 -789 -17 -755
rect 17 -789 33 -755
rect -33 -805 33 -789
rect -30 -836 30 -805
rect -30 -2067 30 -2036
rect -33 -2083 33 -2067
rect -33 -2117 -17 -2083
rect 17 -2117 33 -2083
rect -33 -2133 33 -2117
<< polycont >>
rect -17 2083 17 2117
rect -17 755 17 789
rect -17 647 17 681
rect -17 -681 17 -647
rect -17 -789 17 -755
rect -17 -2117 17 -2083
<< locali >>
rect -190 2185 -94 2219
rect 94 2185 190 2219
rect -190 2123 -156 2185
rect 156 2123 190 2185
rect -33 2083 -17 2117
rect 17 2083 33 2117
rect -76 2024 -42 2040
rect -76 832 -42 848
rect 42 2024 76 2040
rect 42 832 76 848
rect -33 755 -17 789
rect 17 755 33 789
rect -33 647 -17 681
rect 17 647 33 681
rect -76 588 -42 604
rect -76 -604 -42 -588
rect 42 588 76 604
rect 42 -604 76 -588
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -789 -17 -755
rect 17 -789 33 -755
rect -76 -848 -42 -832
rect -76 -2040 -42 -2024
rect 42 -848 76 -832
rect 42 -2040 76 -2024
rect -33 -2117 -17 -2083
rect 17 -2117 33 -2083
rect -190 -2185 -156 -2123
rect 156 -2185 190 -2123
rect -190 -2219 -94 -2185
rect 94 -2219 190 -2185
<< viali >>
rect -17 2083 17 2117
rect -76 848 -42 2024
rect 42 848 76 2024
rect -17 755 17 789
rect -17 647 17 681
rect -76 -588 -42 588
rect 42 -588 76 588
rect -17 -681 17 -647
rect -17 -789 17 -755
rect -76 -2024 -42 -848
rect 42 -2024 76 -848
rect -17 -2117 17 -2083
<< metal1 >>
rect -29 2117 29 2123
rect -29 2083 -17 2117
rect 17 2083 29 2117
rect -29 2077 29 2083
rect -82 2024 -36 2036
rect -82 848 -76 2024
rect -42 848 -36 2024
rect -82 836 -36 848
rect 36 2024 82 2036
rect 36 848 42 2024
rect 76 848 82 2024
rect 36 836 82 848
rect -29 789 29 795
rect -29 755 -17 789
rect 17 755 29 789
rect -29 749 29 755
rect -29 681 29 687
rect -29 647 -17 681
rect 17 647 29 681
rect -29 641 29 647
rect -82 588 -36 600
rect -82 -588 -76 588
rect -42 -588 -36 588
rect -82 -600 -36 -588
rect 36 588 82 600
rect 36 -588 42 588
rect 76 -588 82 588
rect 36 -600 82 -588
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect 17 -681 29 -647
rect -29 -687 29 -681
rect -29 -755 29 -749
rect -29 -789 -17 -755
rect 17 -789 29 -755
rect -29 -795 29 -789
rect -82 -848 -36 -836
rect -82 -2024 -76 -848
rect -42 -2024 -36 -848
rect -82 -2036 -36 -2024
rect 36 -848 82 -836
rect 36 -2024 42 -848
rect 76 -2024 82 -848
rect 36 -2036 82 -2024
rect -29 -2083 29 -2077
rect -29 -2117 -17 -2083
rect 17 -2117 29 -2083
rect -29 -2123 29 -2117
<< properties >>
string FIXED_BBOX -173 -2202 173 2202
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
