magic
tech sky130A
timestamp 1710329453
<< metal1 >>
rect 7205 1812 7305 1912
rect 7205 1612 7305 1712
rect 7205 1412 7305 1512
rect 7205 1212 7305 1312
rect 7205 1012 7305 1112
use pfd  x1
timestamp 1708936645
transform 1 0 5591 0 1 4053
box 393 -940 1978 167
use cp_schem  x2
timestamp 1709641130
transform 1 0 7279 0 1 3524
box 1160 -508 2429 783
use vco  x3
timestamp 1709454227
transform 1 0 8711 0 1 2551
box 1898 -1425 6086 1756
use inverter  x4
timestamp 1709276979
transform 1 0 7766 0 1 3606
box -140 192 520 681
use divider_3N  x5
timestamp 1709895641
transform 1 0 7846 0 1 1610
box 794 -818 2179 205
<< labels >>
flabel metal1 7205 1812 7305 1912 0 FreeSans 128 0 0 0 Ref_sig
port 0 nsew
flabel metal1 7205 1612 7305 1712 0 FreeSans 128 0 0 0 i_bias
port 1 nsew
flabel metal1 7205 1412 7305 1512 0 FreeSans 128 0 0 0 vco_out
port 2 nsew
flabel metal1 7205 1212 7305 1312 0 FreeSans 128 0 0 0 vdd
port 3 nsew
flabel metal1 7205 1012 7305 1112 0 FreeSans 128 0 0 0 vss
port 4 nsew
<< end >>
