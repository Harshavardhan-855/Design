magic
tech sky130A
magscale 1 2
timestamp 1709104634
<< error_p >>
rect -29 2072 29 2078
rect -29 2038 -17 2072
rect -29 2032 29 2038
rect -125 -2038 -67 -2032
rect 67 -2038 125 -2032
rect -125 -2072 -113 -2038
rect 67 -2072 79 -2038
rect -125 -2078 -67 -2072
rect 67 -2078 125 -2072
<< pwell >>
rect -311 -2210 311 2210
<< nmos >>
rect -111 -2000 -81 2000
rect -15 -2000 15 2000
rect 81 -2000 111 2000
<< ndiff >>
rect -173 1988 -111 2000
rect -173 -1988 -161 1988
rect -127 -1988 -111 1988
rect -173 -2000 -111 -1988
rect -81 1988 -15 2000
rect -81 -1988 -65 1988
rect -31 -1988 -15 1988
rect -81 -2000 -15 -1988
rect 15 1988 81 2000
rect 15 -1988 31 1988
rect 65 -1988 81 1988
rect 15 -2000 81 -1988
rect 111 1988 173 2000
rect 111 -1988 127 1988
rect 161 -1988 173 1988
rect 111 -2000 173 -1988
<< ndiffc >>
rect -161 -1988 -127 1988
rect -65 -1988 -31 1988
rect 31 -1988 65 1988
rect 127 -1988 161 1988
<< psubdiff >>
rect -275 2140 -179 2174
rect 179 2140 275 2174
rect -275 2078 -241 2140
rect 241 2078 275 2140
rect -275 -2140 -241 -2078
rect 241 -2140 275 -2078
rect -275 -2174 -179 -2140
rect 179 -2174 275 -2140
<< psubdiffcont >>
rect -179 2140 179 2174
rect -275 -2078 -241 2078
rect 241 -2078 275 2078
rect -179 -2174 179 -2140
<< poly >>
rect -33 2072 33 2088
rect -33 2038 -17 2072
rect 17 2038 33 2072
rect -111 2000 -81 2026
rect -33 2022 33 2038
rect -15 2000 15 2022
rect 81 2000 111 2026
rect -111 -2022 -81 -2000
rect -129 -2038 -63 -2022
rect -15 -2026 15 -2000
rect 81 -2022 111 -2000
rect -129 -2072 -113 -2038
rect -79 -2072 -63 -2038
rect -129 -2088 -63 -2072
rect 63 -2038 129 -2022
rect 63 -2072 79 -2038
rect 113 -2072 129 -2038
rect 63 -2088 129 -2072
<< polycont >>
rect -17 2038 17 2072
rect -113 -2072 -79 -2038
rect 79 -2072 113 -2038
<< locali >>
rect -275 2140 -179 2174
rect 179 2140 275 2174
rect -275 2078 -241 2140
rect 241 2078 275 2140
rect -33 2038 -17 2072
rect 17 2038 33 2072
rect -161 1988 -127 2004
rect -161 -2004 -127 -1988
rect -65 1988 -31 2004
rect -65 -2004 -31 -1988
rect 31 1988 65 2004
rect 31 -2004 65 -1988
rect 127 1988 161 2004
rect 127 -2004 161 -1988
rect -129 -2072 -113 -2038
rect -79 -2072 -63 -2038
rect 63 -2072 79 -2038
rect 113 -2072 129 -2038
rect -275 -2140 -241 -2078
rect 241 -2140 275 -2078
rect -275 -2174 -179 -2140
rect 179 -2174 275 -2140
<< viali >>
rect -17 2038 17 2072
rect -161 -1988 -127 1988
rect -65 -1988 -31 1988
rect 31 -1988 65 1988
rect 127 -1988 161 1988
rect -113 -2072 -79 -2038
rect 79 -2072 113 -2038
<< metal1 >>
rect -29 2072 29 2078
rect -29 2038 -17 2072
rect 17 2038 29 2072
rect -29 2032 29 2038
rect -167 1988 -121 2000
rect -167 -1988 -161 1988
rect -127 -1988 -121 1988
rect -167 -2000 -121 -1988
rect -71 1988 -25 2000
rect -71 -1988 -65 1988
rect -31 -1988 -25 1988
rect -71 -2000 -25 -1988
rect 25 1988 71 2000
rect 25 -1988 31 1988
rect 65 -1988 71 1988
rect 25 -2000 71 -1988
rect 121 1988 167 2000
rect 121 -1988 127 1988
rect 161 -1988 167 1988
rect 121 -2000 167 -1988
rect -125 -2038 -67 -2032
rect -125 -2072 -113 -2038
rect -79 -2072 -67 -2038
rect -125 -2078 -67 -2072
rect 67 -2038 125 -2032
rect 67 -2072 79 -2038
rect 113 -2072 125 -2038
rect 67 -2078 125 -2072
<< properties >>
string FIXED_BBOX -258 -2157 258 2157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
