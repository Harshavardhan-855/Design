* NGSPICE file created from Diffamp.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_po_XJGAA7 a_n100_n680# a_n100_250#
R0 a_n100_250# a_n100_n680# sky130_fd_pr__res_generic_po w=1 l=2.5
.ends

.subckt sky130_fd_pr__nfet_01v8_4H4H2H a_262_n588# a_n328_n588# a_n501_n500# a_561_n500#
+ a_n383_n500# a_498_n588# a_144_n588# a_443_n500# a_n265_n500# a_26_n588# a_n619_n500#
+ a_325_n500# a_n147_n500# a_n210_n588# a_207_n500# a_n564_n588# a_n29_n500# a_n92_n588#
+ a_n721_n674# a_380_n588# a_n446_n588# a_89_n500#
X0 a_n383_n500# a_n446_n588# a_n501_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X1 a_n29_n500# a_n92_n588# a_n147_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X2 a_325_n500# a_262_n588# a_207_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X3 a_n265_n500# a_n328_n588# a_n383_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X4 a_561_n500# a_498_n588# a_443_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.3
X5 a_89_n500# a_26_n588# a_n29_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X6 a_207_n500# a_144_n588# a_89_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X7 a_n501_n500# a_n564_n588# a_n619_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.3
X8 a_n147_n500# a_n210_n588# a_n265_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
X9 a_443_n500# a_380_n588# a_325_n500# a_n721_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.3
.ends

.subckt Diffamp vdd vss inp1 inp2 out2 out1 vbias
XR1 out1 vdd sky130_fd_pr__res_generic_po_XJGAA7
XR2 out2 vdd sky130_fd_pr__res_generic_po_XJGAA7
XXM1 inp1 inp1 m1_n800_604# out1 out1 inp1 inp1 m1_n800_604# m1_n800_604# inp1 out1
+ out1 out1 inp1 m1_n800_604# inp1 m1_n800_604# inp1 vss inp1 inp1 out1 sky130_fd_pr__nfet_01v8_4H4H2H
XXM2 inp2 inp2 m1_n800_604# out2 out2 inp2 inp2 m1_n800_604# m1_n800_604# inp2 out2
+ out2 out2 inp2 m1_n800_604# inp2 m1_n800_604# inp2 vss inp2 inp2 out2 sky130_fd_pr__nfet_01v8_4H4H2H
XXM3 vbias vbias vss m1_n800_604# m1_n800_604# vbias vbias vss vss vbias m1_n800_604#
+ m1_n800_604# m1_n800_604# vbias vss vbias vss vbias vss vbias vbias m1_n800_604#
+ sky130_fd_pr__nfet_01v8_4H4H2H
.ends

