magic
tech sky130A
magscale 1 2
timestamp 1708941600
<< error_p >>
rect -653 144 -595 150
rect -461 144 -403 150
rect -269 144 -211 150
rect -77 144 -19 150
rect 115 144 173 150
rect 307 144 365 150
rect 499 144 557 150
rect 691 144 749 150
rect -653 110 -641 144
rect -461 110 -449 144
rect -269 110 -257 144
rect -77 110 -65 144
rect 115 110 127 144
rect 307 110 319 144
rect 499 110 511 144
rect 691 110 703 144
rect -653 104 -595 110
rect -461 104 -403 110
rect -269 104 -211 110
rect -77 104 -19 110
rect 115 104 173 110
rect 307 104 365 110
rect 499 104 557 110
rect 691 104 749 110
rect -749 -110 -691 -104
rect -557 -110 -499 -104
rect -365 -110 -307 -104
rect -173 -110 -115 -104
rect 19 -110 77 -104
rect 211 -110 269 -104
rect 403 -110 461 -104
rect 595 -110 653 -104
rect -749 -144 -737 -110
rect -557 -144 -545 -110
rect -365 -144 -353 -110
rect -173 -144 -161 -110
rect 19 -144 31 -110
rect 211 -144 223 -110
rect 403 -144 415 -110
rect 595 -144 607 -110
rect -749 -150 -691 -144
rect -557 -150 -499 -144
rect -365 -150 -307 -144
rect -173 -150 -115 -144
rect 19 -150 77 -144
rect 211 -150 269 -144
rect 403 -150 461 -144
rect 595 -150 653 -144
<< nwell >>
rect -935 -282 935 282
<< pmos >>
rect -735 -63 -705 63
rect -639 -63 -609 63
rect -543 -63 -513 63
rect -447 -63 -417 63
rect -351 -63 -321 63
rect -255 -63 -225 63
rect -159 -63 -129 63
rect -63 -63 -33 63
rect 33 -63 63 63
rect 129 -63 159 63
rect 225 -63 255 63
rect 321 -63 351 63
rect 417 -63 447 63
rect 513 -63 543 63
rect 609 -63 639 63
rect 705 -63 735 63
<< pdiff >>
rect -797 51 -735 63
rect -797 -51 -785 51
rect -751 -51 -735 51
rect -797 -63 -735 -51
rect -705 51 -639 63
rect -705 -51 -689 51
rect -655 -51 -639 51
rect -705 -63 -639 -51
rect -609 51 -543 63
rect -609 -51 -593 51
rect -559 -51 -543 51
rect -609 -63 -543 -51
rect -513 51 -447 63
rect -513 -51 -497 51
rect -463 -51 -447 51
rect -513 -63 -447 -51
rect -417 51 -351 63
rect -417 -51 -401 51
rect -367 -51 -351 51
rect -417 -63 -351 -51
rect -321 51 -255 63
rect -321 -51 -305 51
rect -271 -51 -255 51
rect -321 -63 -255 -51
rect -225 51 -159 63
rect -225 -51 -209 51
rect -175 -51 -159 51
rect -225 -63 -159 -51
rect -129 51 -63 63
rect -129 -51 -113 51
rect -79 -51 -63 51
rect -129 -63 -63 -51
rect -33 51 33 63
rect -33 -51 -17 51
rect 17 -51 33 51
rect -33 -63 33 -51
rect 63 51 129 63
rect 63 -51 79 51
rect 113 -51 129 51
rect 63 -63 129 -51
rect 159 51 225 63
rect 159 -51 175 51
rect 209 -51 225 51
rect 159 -63 225 -51
rect 255 51 321 63
rect 255 -51 271 51
rect 305 -51 321 51
rect 255 -63 321 -51
rect 351 51 417 63
rect 351 -51 367 51
rect 401 -51 417 51
rect 351 -63 417 -51
rect 447 51 513 63
rect 447 -51 463 51
rect 497 -51 513 51
rect 447 -63 513 -51
rect 543 51 609 63
rect 543 -51 559 51
rect 593 -51 609 51
rect 543 -63 609 -51
rect 639 51 705 63
rect 639 -51 655 51
rect 689 -51 705 51
rect 639 -63 705 -51
rect 735 51 797 63
rect 735 -51 751 51
rect 785 -51 797 51
rect 735 -63 797 -51
<< pdiffc >>
rect -785 -51 -751 51
rect -689 -51 -655 51
rect -593 -51 -559 51
rect -497 -51 -463 51
rect -401 -51 -367 51
rect -305 -51 -271 51
rect -209 -51 -175 51
rect -113 -51 -79 51
rect -17 -51 17 51
rect 79 -51 113 51
rect 175 -51 209 51
rect 271 -51 305 51
rect 367 -51 401 51
rect 463 -51 497 51
rect 559 -51 593 51
rect 655 -51 689 51
rect 751 -51 785 51
<< nsubdiff >>
rect -899 212 -803 246
rect 803 212 899 246
rect -899 150 -865 212
rect 865 150 899 212
rect -899 -212 -865 -150
rect 865 -212 899 -150
rect -899 -246 -803 -212
rect 803 -246 899 -212
<< nsubdiffcont >>
rect -803 212 803 246
rect -899 -150 -865 150
rect 865 -150 899 150
rect -803 -246 803 -212
<< poly >>
rect -657 144 -591 160
rect -657 110 -641 144
rect -607 110 -591 144
rect -657 94 -591 110
rect -465 144 -399 160
rect -465 110 -449 144
rect -415 110 -399 144
rect -465 94 -399 110
rect -273 144 -207 160
rect -273 110 -257 144
rect -223 110 -207 144
rect -273 94 -207 110
rect -81 144 -15 160
rect -81 110 -65 144
rect -31 110 -15 144
rect -81 94 -15 110
rect 111 144 177 160
rect 111 110 127 144
rect 161 110 177 144
rect 111 94 177 110
rect 303 144 369 160
rect 303 110 319 144
rect 353 110 369 144
rect 303 94 369 110
rect 495 144 561 160
rect 495 110 511 144
rect 545 110 561 144
rect 495 94 561 110
rect 687 144 753 160
rect 687 110 703 144
rect 737 110 753 144
rect 687 94 753 110
rect -735 63 -705 89
rect -639 63 -609 94
rect -543 63 -513 89
rect -447 63 -417 94
rect -351 63 -321 89
rect -255 63 -225 94
rect -159 63 -129 89
rect -63 63 -33 94
rect 33 63 63 89
rect 129 63 159 94
rect 225 63 255 89
rect 321 63 351 94
rect 417 63 447 89
rect 513 63 543 94
rect 609 63 639 89
rect 705 63 735 94
rect -735 -94 -705 -63
rect -639 -89 -609 -63
rect -543 -94 -513 -63
rect -447 -89 -417 -63
rect -351 -94 -321 -63
rect -255 -89 -225 -63
rect -159 -94 -129 -63
rect -63 -89 -33 -63
rect 33 -94 63 -63
rect 129 -89 159 -63
rect 225 -94 255 -63
rect 321 -89 351 -63
rect 417 -94 447 -63
rect 513 -89 543 -63
rect 609 -94 639 -63
rect 705 -89 735 -63
rect -753 -110 -687 -94
rect -753 -144 -737 -110
rect -703 -144 -687 -110
rect -753 -160 -687 -144
rect -561 -110 -495 -94
rect -561 -144 -545 -110
rect -511 -144 -495 -110
rect -561 -160 -495 -144
rect -369 -110 -303 -94
rect -369 -144 -353 -110
rect -319 -144 -303 -110
rect -369 -160 -303 -144
rect -177 -110 -111 -94
rect -177 -144 -161 -110
rect -127 -144 -111 -110
rect -177 -160 -111 -144
rect 15 -110 81 -94
rect 15 -144 31 -110
rect 65 -144 81 -110
rect 15 -160 81 -144
rect 207 -110 273 -94
rect 207 -144 223 -110
rect 257 -144 273 -110
rect 207 -160 273 -144
rect 399 -110 465 -94
rect 399 -144 415 -110
rect 449 -144 465 -110
rect 399 -160 465 -144
rect 591 -110 657 -94
rect 591 -144 607 -110
rect 641 -144 657 -110
rect 591 -160 657 -144
<< polycont >>
rect -641 110 -607 144
rect -449 110 -415 144
rect -257 110 -223 144
rect -65 110 -31 144
rect 127 110 161 144
rect 319 110 353 144
rect 511 110 545 144
rect 703 110 737 144
rect -737 -144 -703 -110
rect -545 -144 -511 -110
rect -353 -144 -319 -110
rect -161 -144 -127 -110
rect 31 -144 65 -110
rect 223 -144 257 -110
rect 415 -144 449 -110
rect 607 -144 641 -110
<< locali >>
rect -899 212 -803 246
rect 803 212 899 246
rect -899 150 -865 212
rect 865 150 899 212
rect -657 110 -641 144
rect -607 110 -591 144
rect -465 110 -449 144
rect -415 110 -399 144
rect -273 110 -257 144
rect -223 110 -207 144
rect -81 110 -65 144
rect -31 110 -15 144
rect 111 110 127 144
rect 161 110 177 144
rect 303 110 319 144
rect 353 110 369 144
rect 495 110 511 144
rect 545 110 561 144
rect 687 110 703 144
rect 737 110 753 144
rect -785 51 -751 67
rect -785 -67 -751 -51
rect -689 51 -655 67
rect -689 -67 -655 -51
rect -593 51 -559 67
rect -593 -67 -559 -51
rect -497 51 -463 67
rect -497 -67 -463 -51
rect -401 51 -367 67
rect -401 -67 -367 -51
rect -305 51 -271 67
rect -305 -67 -271 -51
rect -209 51 -175 67
rect -209 -67 -175 -51
rect -113 51 -79 67
rect -113 -67 -79 -51
rect -17 51 17 67
rect -17 -67 17 -51
rect 79 51 113 67
rect 79 -67 113 -51
rect 175 51 209 67
rect 175 -67 209 -51
rect 271 51 305 67
rect 271 -67 305 -51
rect 367 51 401 67
rect 367 -67 401 -51
rect 463 51 497 67
rect 463 -67 497 -51
rect 559 51 593 67
rect 559 -67 593 -51
rect 655 51 689 67
rect 655 -67 689 -51
rect 751 51 785 67
rect 751 -67 785 -51
rect -753 -144 -737 -110
rect -703 -144 -687 -110
rect -561 -144 -545 -110
rect -511 -144 -495 -110
rect -369 -144 -353 -110
rect -319 -144 -303 -110
rect -177 -144 -161 -110
rect -127 -144 -111 -110
rect 15 -144 31 -110
rect 65 -144 81 -110
rect 207 -144 223 -110
rect 257 -144 273 -110
rect 399 -144 415 -110
rect 449 -144 465 -110
rect 591 -144 607 -110
rect 641 -144 657 -110
rect -899 -212 -865 -150
rect 865 -212 899 -150
rect -899 -246 -803 -212
rect 803 -246 899 -212
<< viali >>
rect -641 110 -607 144
rect -449 110 -415 144
rect -257 110 -223 144
rect -65 110 -31 144
rect 127 110 161 144
rect 319 110 353 144
rect 511 110 545 144
rect 703 110 737 144
rect -785 -51 -751 51
rect -689 -51 -655 51
rect -593 -51 -559 51
rect -497 -51 -463 51
rect -401 -51 -367 51
rect -305 -51 -271 51
rect -209 -51 -175 51
rect -113 -51 -79 51
rect -17 -51 17 51
rect 79 -51 113 51
rect 175 -51 209 51
rect 271 -51 305 51
rect 367 -51 401 51
rect 463 -51 497 51
rect 559 -51 593 51
rect 655 -51 689 51
rect 751 -51 785 51
rect -737 -144 -703 -110
rect -545 -144 -511 -110
rect -353 -144 -319 -110
rect -161 -144 -127 -110
rect 31 -144 65 -110
rect 223 -144 257 -110
rect 415 -144 449 -110
rect 607 -144 641 -110
<< metal1 >>
rect -653 144 -595 150
rect -653 110 -641 144
rect -607 110 -595 144
rect -653 104 -595 110
rect -461 144 -403 150
rect -461 110 -449 144
rect -415 110 -403 144
rect -461 104 -403 110
rect -269 144 -211 150
rect -269 110 -257 144
rect -223 110 -211 144
rect -269 104 -211 110
rect -77 144 -19 150
rect -77 110 -65 144
rect -31 110 -19 144
rect -77 104 -19 110
rect 115 144 173 150
rect 115 110 127 144
rect 161 110 173 144
rect 115 104 173 110
rect 307 144 365 150
rect 307 110 319 144
rect 353 110 365 144
rect 307 104 365 110
rect 499 144 557 150
rect 499 110 511 144
rect 545 110 557 144
rect 499 104 557 110
rect 691 144 749 150
rect 691 110 703 144
rect 737 110 749 144
rect 691 104 749 110
rect -791 51 -745 63
rect -791 -51 -785 51
rect -751 -51 -745 51
rect -791 -63 -745 -51
rect -695 51 -649 63
rect -695 -51 -689 51
rect -655 -51 -649 51
rect -695 -63 -649 -51
rect -599 51 -553 63
rect -599 -51 -593 51
rect -559 -51 -553 51
rect -599 -63 -553 -51
rect -503 51 -457 63
rect -503 -51 -497 51
rect -463 -51 -457 51
rect -503 -63 -457 -51
rect -407 51 -361 63
rect -407 -51 -401 51
rect -367 -51 -361 51
rect -407 -63 -361 -51
rect -311 51 -265 63
rect -311 -51 -305 51
rect -271 -51 -265 51
rect -311 -63 -265 -51
rect -215 51 -169 63
rect -215 -51 -209 51
rect -175 -51 -169 51
rect -215 -63 -169 -51
rect -119 51 -73 63
rect -119 -51 -113 51
rect -79 -51 -73 51
rect -119 -63 -73 -51
rect -23 51 23 63
rect -23 -51 -17 51
rect 17 -51 23 51
rect -23 -63 23 -51
rect 73 51 119 63
rect 73 -51 79 51
rect 113 -51 119 51
rect 73 -63 119 -51
rect 169 51 215 63
rect 169 -51 175 51
rect 209 -51 215 51
rect 169 -63 215 -51
rect 265 51 311 63
rect 265 -51 271 51
rect 305 -51 311 51
rect 265 -63 311 -51
rect 361 51 407 63
rect 361 -51 367 51
rect 401 -51 407 51
rect 361 -63 407 -51
rect 457 51 503 63
rect 457 -51 463 51
rect 497 -51 503 51
rect 457 -63 503 -51
rect 553 51 599 63
rect 553 -51 559 51
rect 593 -51 599 51
rect 553 -63 599 -51
rect 649 51 695 63
rect 649 -51 655 51
rect 689 -51 695 51
rect 649 -63 695 -51
rect 745 51 791 63
rect 745 -51 751 51
rect 785 -51 791 51
rect 745 -63 791 -51
rect -749 -110 -691 -104
rect -749 -144 -737 -110
rect -703 -144 -691 -110
rect -749 -150 -691 -144
rect -557 -110 -499 -104
rect -557 -144 -545 -110
rect -511 -144 -499 -110
rect -557 -150 -499 -144
rect -365 -110 -307 -104
rect -365 -144 -353 -110
rect -319 -144 -307 -110
rect -365 -150 -307 -144
rect -173 -110 -115 -104
rect -173 -144 -161 -110
rect -127 -144 -115 -110
rect -173 -150 -115 -144
rect 19 -110 77 -104
rect 19 -144 31 -110
rect 65 -144 77 -110
rect 19 -150 77 -144
rect 211 -110 269 -104
rect 211 -144 223 -110
rect 257 -144 269 -110
rect 211 -150 269 -144
rect 403 -110 461 -104
rect 403 -144 415 -110
rect 449 -144 461 -110
rect 403 -150 461 -144
rect 595 -110 653 -104
rect 595 -144 607 -110
rect 641 -144 653 -110
rect 595 -150 653 -144
<< properties >>
string FIXED_BBOX -882 -229 882 229
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.625 l 0.15 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
