magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -365 171 -307 177
rect -173 171 -115 177
rect 19 171 77 177
rect 211 171 269 177
rect 403 171 461 177
rect -365 137 -353 171
rect -173 137 -161 171
rect 19 137 31 171
rect 211 137 223 171
rect 403 137 415 171
rect -365 131 -307 137
rect -173 131 -115 137
rect 19 131 77 137
rect 211 131 269 137
rect 403 131 461 137
rect -461 -137 -403 -131
rect -269 -137 -211 -131
rect -77 -137 -19 -131
rect 115 -137 173 -131
rect 307 -137 365 -131
rect -461 -171 -449 -137
rect -269 -171 -257 -137
rect -77 -171 -65 -137
rect 115 -171 127 -137
rect 307 -171 319 -137
rect -461 -177 -403 -171
rect -269 -177 -211 -171
rect -77 -177 -19 -171
rect 115 -177 173 -171
rect 307 -177 365 -171
<< nwell >>
rect -647 -309 647 309
<< pmos >>
rect -447 -90 -417 90
rect -351 -90 -321 90
rect -255 -90 -225 90
rect -159 -90 -129 90
rect -63 -90 -33 90
rect 33 -90 63 90
rect 129 -90 159 90
rect 225 -90 255 90
rect 321 -90 351 90
rect 417 -90 447 90
<< pdiff >>
rect -509 78 -447 90
rect -509 -78 -497 78
rect -463 -78 -447 78
rect -509 -90 -447 -78
rect -417 78 -351 90
rect -417 -78 -401 78
rect -367 -78 -351 78
rect -417 -90 -351 -78
rect -321 78 -255 90
rect -321 -78 -305 78
rect -271 -78 -255 78
rect -321 -90 -255 -78
rect -225 78 -159 90
rect -225 -78 -209 78
rect -175 -78 -159 78
rect -225 -90 -159 -78
rect -129 78 -63 90
rect -129 -78 -113 78
rect -79 -78 -63 78
rect -129 -90 -63 -78
rect -33 78 33 90
rect -33 -78 -17 78
rect 17 -78 33 78
rect -33 -90 33 -78
rect 63 78 129 90
rect 63 -78 79 78
rect 113 -78 129 78
rect 63 -90 129 -78
rect 159 78 225 90
rect 159 -78 175 78
rect 209 -78 225 78
rect 159 -90 225 -78
rect 255 78 321 90
rect 255 -78 271 78
rect 305 -78 321 78
rect 255 -90 321 -78
rect 351 78 417 90
rect 351 -78 367 78
rect 401 -78 417 78
rect 351 -90 417 -78
rect 447 78 509 90
rect 447 -78 463 78
rect 497 -78 509 78
rect 447 -90 509 -78
<< pdiffc >>
rect -497 -78 -463 78
rect -401 -78 -367 78
rect -305 -78 -271 78
rect -209 -78 -175 78
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
rect 175 -78 209 78
rect 271 -78 305 78
rect 367 -78 401 78
rect 463 -78 497 78
<< nsubdiff >>
rect -611 239 -515 273
rect 515 239 611 273
rect -611 177 -577 239
rect 577 177 611 239
rect -611 -239 -577 -177
rect 577 -239 611 -177
rect -611 -273 -515 -239
rect 515 -273 611 -239
<< nsubdiffcont >>
rect -515 239 515 273
rect -611 -177 -577 177
rect 577 -177 611 177
rect -515 -273 515 -239
<< poly >>
rect -369 171 -303 187
rect -369 137 -353 171
rect -319 137 -303 171
rect -369 121 -303 137
rect -177 171 -111 187
rect -177 137 -161 171
rect -127 137 -111 171
rect -177 121 -111 137
rect 15 171 81 187
rect 15 137 31 171
rect 65 137 81 171
rect 15 121 81 137
rect 207 171 273 187
rect 207 137 223 171
rect 257 137 273 171
rect 207 121 273 137
rect 399 171 465 187
rect 399 137 415 171
rect 449 137 465 171
rect 399 121 465 137
rect -447 90 -417 116
rect -351 90 -321 121
rect -255 90 -225 116
rect -159 90 -129 121
rect -63 90 -33 116
rect 33 90 63 121
rect 129 90 159 116
rect 225 90 255 121
rect 321 90 351 116
rect 417 90 447 121
rect -447 -121 -417 -90
rect -351 -116 -321 -90
rect -255 -121 -225 -90
rect -159 -116 -129 -90
rect -63 -121 -33 -90
rect 33 -116 63 -90
rect 129 -121 159 -90
rect 225 -116 255 -90
rect 321 -121 351 -90
rect 417 -116 447 -90
rect -465 -137 -399 -121
rect -465 -171 -449 -137
rect -415 -171 -399 -137
rect -465 -187 -399 -171
rect -273 -137 -207 -121
rect -273 -171 -257 -137
rect -223 -171 -207 -137
rect -273 -187 -207 -171
rect -81 -137 -15 -121
rect -81 -171 -65 -137
rect -31 -171 -15 -137
rect -81 -187 -15 -171
rect 111 -137 177 -121
rect 111 -171 127 -137
rect 161 -171 177 -137
rect 111 -187 177 -171
rect 303 -137 369 -121
rect 303 -171 319 -137
rect 353 -171 369 -137
rect 303 -187 369 -171
<< polycont >>
rect -353 137 -319 171
rect -161 137 -127 171
rect 31 137 65 171
rect 223 137 257 171
rect 415 137 449 171
rect -449 -171 -415 -137
rect -257 -171 -223 -137
rect -65 -171 -31 -137
rect 127 -171 161 -137
rect 319 -171 353 -137
<< locali >>
rect -611 239 -515 273
rect 515 239 611 273
rect -611 177 -577 239
rect 577 177 611 239
rect -369 137 -353 171
rect -319 137 -303 171
rect -177 137 -161 171
rect -127 137 -111 171
rect 15 137 31 171
rect 65 137 81 171
rect 207 137 223 171
rect 257 137 273 171
rect 399 137 415 171
rect 449 137 465 171
rect -497 78 -463 94
rect -497 -94 -463 -78
rect -401 78 -367 94
rect -401 -94 -367 -78
rect -305 78 -271 94
rect -305 -94 -271 -78
rect -209 78 -175 94
rect -209 -94 -175 -78
rect -113 78 -79 94
rect -113 -94 -79 -78
rect -17 78 17 94
rect -17 -94 17 -78
rect 79 78 113 94
rect 79 -94 113 -78
rect 175 78 209 94
rect 175 -94 209 -78
rect 271 78 305 94
rect 271 -94 305 -78
rect 367 78 401 94
rect 367 -94 401 -78
rect 463 78 497 94
rect 463 -94 497 -78
rect -465 -171 -449 -137
rect -415 -171 -399 -137
rect -273 -171 -257 -137
rect -223 -171 -207 -137
rect -81 -171 -65 -137
rect -31 -171 -15 -137
rect 111 -171 127 -137
rect 161 -171 177 -137
rect 303 -171 319 -137
rect 353 -171 369 -137
rect -611 -239 -577 -177
rect 577 -239 611 -177
rect -611 -273 -515 -239
rect 515 -273 611 -239
<< viali >>
rect -353 137 -319 171
rect -161 137 -127 171
rect 31 137 65 171
rect 223 137 257 171
rect 415 137 449 171
rect -497 -78 -463 78
rect -401 -78 -367 78
rect -305 -78 -271 78
rect -209 -78 -175 78
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
rect 175 -78 209 78
rect 271 -78 305 78
rect 367 -78 401 78
rect 463 -78 497 78
rect -449 -171 -415 -137
rect -257 -171 -223 -137
rect -65 -171 -31 -137
rect 127 -171 161 -137
rect 319 -171 353 -137
<< metal1 >>
rect -365 171 -307 177
rect -365 137 -353 171
rect -319 137 -307 171
rect -365 131 -307 137
rect -173 171 -115 177
rect -173 137 -161 171
rect -127 137 -115 171
rect -173 131 -115 137
rect 19 171 77 177
rect 19 137 31 171
rect 65 137 77 171
rect 19 131 77 137
rect 211 171 269 177
rect 211 137 223 171
rect 257 137 269 171
rect 211 131 269 137
rect 403 171 461 177
rect 403 137 415 171
rect 449 137 461 171
rect 403 131 461 137
rect -503 78 -457 90
rect -503 -78 -497 78
rect -463 -78 -457 78
rect -503 -90 -457 -78
rect -407 78 -361 90
rect -407 -78 -401 78
rect -367 -78 -361 78
rect -407 -90 -361 -78
rect -311 78 -265 90
rect -311 -78 -305 78
rect -271 -78 -265 78
rect -311 -90 -265 -78
rect -215 78 -169 90
rect -215 -78 -209 78
rect -175 -78 -169 78
rect -215 -90 -169 -78
rect -119 78 -73 90
rect -119 -78 -113 78
rect -79 -78 -73 78
rect -119 -90 -73 -78
rect -23 78 23 90
rect -23 -78 -17 78
rect 17 -78 23 78
rect -23 -90 23 -78
rect 73 78 119 90
rect 73 -78 79 78
rect 113 -78 119 78
rect 73 -90 119 -78
rect 169 78 215 90
rect 169 -78 175 78
rect 209 -78 215 78
rect 169 -90 215 -78
rect 265 78 311 90
rect 265 -78 271 78
rect 305 -78 311 78
rect 265 -90 311 -78
rect 361 78 407 90
rect 361 -78 367 78
rect 401 -78 407 78
rect 361 -90 407 -78
rect 457 78 503 90
rect 457 -78 463 78
rect 497 -78 503 78
rect 457 -90 503 -78
rect -461 -137 -403 -131
rect -461 -171 -449 -137
rect -415 -171 -403 -137
rect -461 -177 -403 -171
rect -269 -137 -211 -131
rect -269 -171 -257 -137
rect -223 -171 -211 -137
rect -269 -177 -211 -171
rect -77 -137 -19 -131
rect -77 -171 -65 -137
rect -31 -171 -19 -137
rect -77 -177 -19 -171
rect 115 -137 173 -131
rect 115 -171 127 -137
rect 161 -171 173 -137
rect 115 -177 173 -171
rect 307 -137 365 -131
rect 307 -171 319 -137
rect 353 -171 365 -137
rect 307 -177 365 -171
<< properties >>
string FIXED_BBOX -594 -256 594 256
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.9 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
