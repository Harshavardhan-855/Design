magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< pwell >>
rect -1057 -360 1057 360
<< nmos >>
rect -861 -150 -741 150
rect -683 -150 -563 150
rect -505 -150 -385 150
rect -327 -150 -207 150
rect -149 -150 -29 150
rect 29 -150 149 150
rect 207 -150 327 150
rect 385 -150 505 150
rect 563 -150 683 150
rect 741 -150 861 150
<< ndiff >>
rect -919 138 -861 150
rect -919 -138 -907 138
rect -873 -138 -861 138
rect -919 -150 -861 -138
rect -741 138 -683 150
rect -741 -138 -729 138
rect -695 -138 -683 138
rect -741 -150 -683 -138
rect -563 138 -505 150
rect -563 -138 -551 138
rect -517 -138 -505 138
rect -563 -150 -505 -138
rect -385 138 -327 150
rect -385 -138 -373 138
rect -339 -138 -327 138
rect -385 -150 -327 -138
rect -207 138 -149 150
rect -207 -138 -195 138
rect -161 -138 -149 138
rect -207 -150 -149 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 149 138 207 150
rect 149 -138 161 138
rect 195 -138 207 138
rect 149 -150 207 -138
rect 327 138 385 150
rect 327 -138 339 138
rect 373 -138 385 138
rect 327 -150 385 -138
rect 505 138 563 150
rect 505 -138 517 138
rect 551 -138 563 138
rect 505 -150 563 -138
rect 683 138 741 150
rect 683 -138 695 138
rect 729 -138 741 138
rect 683 -150 741 -138
rect 861 138 919 150
rect 861 -138 873 138
rect 907 -138 919 138
rect 861 -150 919 -138
<< ndiffc >>
rect -907 -138 -873 138
rect -729 -138 -695 138
rect -551 -138 -517 138
rect -373 -138 -339 138
rect -195 -138 -161 138
rect -17 -138 17 138
rect 161 -138 195 138
rect 339 -138 373 138
rect 517 -138 551 138
rect 695 -138 729 138
rect 873 -138 907 138
<< psubdiff >>
rect -1021 290 -925 324
rect 925 290 1021 324
rect -1021 228 -987 290
rect 987 228 1021 290
rect -1021 -290 -987 -228
rect 987 -290 1021 -228
rect -1021 -324 -925 -290
rect 925 -324 1021 -290
<< psubdiffcont >>
rect -925 290 925 324
rect -1021 -228 -987 228
rect 987 -228 1021 228
rect -925 -324 925 -290
<< poly >>
rect -861 222 -741 238
rect -861 188 -845 222
rect -757 188 -741 222
rect -861 150 -741 188
rect -683 222 -563 238
rect -683 188 -667 222
rect -579 188 -563 222
rect -683 150 -563 188
rect -505 222 -385 238
rect -505 188 -489 222
rect -401 188 -385 222
rect -505 150 -385 188
rect -327 222 -207 238
rect -327 188 -311 222
rect -223 188 -207 222
rect -327 150 -207 188
rect -149 222 -29 238
rect -149 188 -133 222
rect -45 188 -29 222
rect -149 150 -29 188
rect 29 222 149 238
rect 29 188 45 222
rect 133 188 149 222
rect 29 150 149 188
rect 207 222 327 238
rect 207 188 223 222
rect 311 188 327 222
rect 207 150 327 188
rect 385 222 505 238
rect 385 188 401 222
rect 489 188 505 222
rect 385 150 505 188
rect 563 222 683 238
rect 563 188 579 222
rect 667 188 683 222
rect 563 150 683 188
rect 741 222 861 238
rect 741 188 757 222
rect 845 188 861 222
rect 741 150 861 188
rect -861 -188 -741 -150
rect -861 -222 -845 -188
rect -757 -222 -741 -188
rect -861 -238 -741 -222
rect -683 -188 -563 -150
rect -683 -222 -667 -188
rect -579 -222 -563 -188
rect -683 -238 -563 -222
rect -505 -188 -385 -150
rect -505 -222 -489 -188
rect -401 -222 -385 -188
rect -505 -238 -385 -222
rect -327 -188 -207 -150
rect -327 -222 -311 -188
rect -223 -222 -207 -188
rect -327 -238 -207 -222
rect -149 -188 -29 -150
rect -149 -222 -133 -188
rect -45 -222 -29 -188
rect -149 -238 -29 -222
rect 29 -188 149 -150
rect 29 -222 45 -188
rect 133 -222 149 -188
rect 29 -238 149 -222
rect 207 -188 327 -150
rect 207 -222 223 -188
rect 311 -222 327 -188
rect 207 -238 327 -222
rect 385 -188 505 -150
rect 385 -222 401 -188
rect 489 -222 505 -188
rect 385 -238 505 -222
rect 563 -188 683 -150
rect 563 -222 579 -188
rect 667 -222 683 -188
rect 563 -238 683 -222
rect 741 -188 861 -150
rect 741 -222 757 -188
rect 845 -222 861 -188
rect 741 -238 861 -222
<< polycont >>
rect -845 188 -757 222
rect -667 188 -579 222
rect -489 188 -401 222
rect -311 188 -223 222
rect -133 188 -45 222
rect 45 188 133 222
rect 223 188 311 222
rect 401 188 489 222
rect 579 188 667 222
rect 757 188 845 222
rect -845 -222 -757 -188
rect -667 -222 -579 -188
rect -489 -222 -401 -188
rect -311 -222 -223 -188
rect -133 -222 -45 -188
rect 45 -222 133 -188
rect 223 -222 311 -188
rect 401 -222 489 -188
rect 579 -222 667 -188
rect 757 -222 845 -188
<< locali >>
rect -1021 290 -925 324
rect 925 290 1021 324
rect -1021 228 -987 290
rect 987 228 1021 290
rect -861 188 -845 222
rect -757 188 -741 222
rect -683 188 -667 222
rect -579 188 -563 222
rect -505 188 -489 222
rect -401 188 -385 222
rect -327 188 -311 222
rect -223 188 -207 222
rect -149 188 -133 222
rect -45 188 -29 222
rect 29 188 45 222
rect 133 188 149 222
rect 207 188 223 222
rect 311 188 327 222
rect 385 188 401 222
rect 489 188 505 222
rect 563 188 579 222
rect 667 188 683 222
rect 741 188 757 222
rect 845 188 861 222
rect -907 138 -873 154
rect -907 -154 -873 -138
rect -729 138 -695 154
rect -729 -154 -695 -138
rect -551 138 -517 154
rect -551 -154 -517 -138
rect -373 138 -339 154
rect -373 -154 -339 -138
rect -195 138 -161 154
rect -195 -154 -161 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 161 138 195 154
rect 161 -154 195 -138
rect 339 138 373 154
rect 339 -154 373 -138
rect 517 138 551 154
rect 517 -154 551 -138
rect 695 138 729 154
rect 695 -154 729 -138
rect 873 138 907 154
rect 873 -154 907 -138
rect -861 -222 -845 -188
rect -757 -222 -741 -188
rect -683 -222 -667 -188
rect -579 -222 -563 -188
rect -505 -222 -489 -188
rect -401 -222 -385 -188
rect -327 -222 -311 -188
rect -223 -222 -207 -188
rect -149 -222 -133 -188
rect -45 -222 -29 -188
rect 29 -222 45 -188
rect 133 -222 149 -188
rect 207 -222 223 -188
rect 311 -222 327 -188
rect 385 -222 401 -188
rect 489 -222 505 -188
rect 563 -222 579 -188
rect 667 -222 683 -188
rect 741 -222 757 -188
rect 845 -222 861 -188
rect -1021 -290 -987 -228
rect 987 -290 1021 -228
rect -1021 -324 -925 -290
rect 925 -324 1021 -290
<< viali >>
rect -845 188 -757 222
rect -667 188 -579 222
rect -489 188 -401 222
rect -311 188 -223 222
rect -133 188 -45 222
rect 45 188 133 222
rect 223 188 311 222
rect 401 188 489 222
rect 579 188 667 222
rect 757 188 845 222
rect -907 -138 -873 138
rect -729 -138 -695 138
rect -551 -138 -517 138
rect -373 -138 -339 138
rect -195 -138 -161 138
rect -17 -138 17 138
rect 161 -138 195 138
rect 339 -138 373 138
rect 517 -138 551 138
rect 695 -138 729 138
rect 873 -138 907 138
rect -845 -222 -757 -188
rect -667 -222 -579 -188
rect -489 -222 -401 -188
rect -311 -222 -223 -188
rect -133 -222 -45 -188
rect 45 -222 133 -188
rect 223 -222 311 -188
rect 401 -222 489 -188
rect 579 -222 667 -188
rect 757 -222 845 -188
<< metal1 >>
rect -857 222 -745 228
rect -857 188 -845 222
rect -757 188 -745 222
rect -857 182 -745 188
rect -679 222 -567 228
rect -679 188 -667 222
rect -579 188 -567 222
rect -679 182 -567 188
rect -501 222 -389 228
rect -501 188 -489 222
rect -401 188 -389 222
rect -501 182 -389 188
rect -323 222 -211 228
rect -323 188 -311 222
rect -223 188 -211 222
rect -323 182 -211 188
rect -145 222 -33 228
rect -145 188 -133 222
rect -45 188 -33 222
rect -145 182 -33 188
rect 33 222 145 228
rect 33 188 45 222
rect 133 188 145 222
rect 33 182 145 188
rect 211 222 323 228
rect 211 188 223 222
rect 311 188 323 222
rect 211 182 323 188
rect 389 222 501 228
rect 389 188 401 222
rect 489 188 501 222
rect 389 182 501 188
rect 567 222 679 228
rect 567 188 579 222
rect 667 188 679 222
rect 567 182 679 188
rect 745 222 857 228
rect 745 188 757 222
rect 845 188 857 222
rect 745 182 857 188
rect -913 138 -867 150
rect -913 -138 -907 138
rect -873 -138 -867 138
rect -913 -150 -867 -138
rect -735 138 -689 150
rect -735 -138 -729 138
rect -695 -138 -689 138
rect -735 -150 -689 -138
rect -557 138 -511 150
rect -557 -138 -551 138
rect -517 -138 -511 138
rect -557 -150 -511 -138
rect -379 138 -333 150
rect -379 -138 -373 138
rect -339 -138 -333 138
rect -379 -150 -333 -138
rect -201 138 -155 150
rect -201 -138 -195 138
rect -161 -138 -155 138
rect -201 -150 -155 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 155 138 201 150
rect 155 -138 161 138
rect 195 -138 201 138
rect 155 -150 201 -138
rect 333 138 379 150
rect 333 -138 339 138
rect 373 -138 379 138
rect 333 -150 379 -138
rect 511 138 557 150
rect 511 -138 517 138
rect 551 -138 557 138
rect 511 -150 557 -138
rect 689 138 735 150
rect 689 -138 695 138
rect 729 -138 735 138
rect 689 -150 735 -138
rect 867 138 913 150
rect 867 -138 873 138
rect 907 -138 913 138
rect 867 -150 913 -138
rect -857 -188 -745 -182
rect -857 -222 -845 -188
rect -757 -222 -745 -188
rect -857 -228 -745 -222
rect -679 -188 -567 -182
rect -679 -222 -667 -188
rect -579 -222 -567 -188
rect -679 -228 -567 -222
rect -501 -188 -389 -182
rect -501 -222 -489 -188
rect -401 -222 -389 -188
rect -501 -228 -389 -222
rect -323 -188 -211 -182
rect -323 -222 -311 -188
rect -223 -222 -211 -188
rect -323 -228 -211 -222
rect -145 -188 -33 -182
rect -145 -222 -133 -188
rect -45 -222 -33 -188
rect -145 -228 -33 -222
rect 33 -188 145 -182
rect 33 -222 45 -188
rect 133 -222 145 -188
rect 33 -228 145 -222
rect 211 -188 323 -182
rect 211 -222 223 -188
rect 311 -222 323 -188
rect 211 -228 323 -222
rect 389 -188 501 -182
rect 389 -222 401 -188
rect 489 -222 501 -188
rect 389 -228 501 -222
rect 567 -188 679 -182
rect 567 -222 579 -188
rect 667 -222 679 -188
rect 567 -228 679 -222
rect 745 -188 857 -182
rect 745 -222 757 -188
rect 845 -222 857 -188
rect 745 -228 857 -222
<< properties >>
string FIXED_BBOX -1004 -307 1004 307
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.5 l 0.6 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
