magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< pwell >>
rect -1057 -252 1057 252
<< nmos >>
rect -861 -42 -741 42
rect -683 -42 -563 42
rect -505 -42 -385 42
rect -327 -42 -207 42
rect -149 -42 -29 42
rect 29 -42 149 42
rect 207 -42 327 42
rect 385 -42 505 42
rect 563 -42 683 42
rect 741 -42 861 42
<< ndiff >>
rect -919 30 -861 42
rect -919 -30 -907 30
rect -873 -30 -861 30
rect -919 -42 -861 -30
rect -741 30 -683 42
rect -741 -30 -729 30
rect -695 -30 -683 30
rect -741 -42 -683 -30
rect -563 30 -505 42
rect -563 -30 -551 30
rect -517 -30 -505 30
rect -563 -42 -505 -30
rect -385 30 -327 42
rect -385 -30 -373 30
rect -339 -30 -327 30
rect -385 -42 -327 -30
rect -207 30 -149 42
rect -207 -30 -195 30
rect -161 -30 -149 30
rect -207 -42 -149 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 149 30 207 42
rect 149 -30 161 30
rect 195 -30 207 30
rect 149 -42 207 -30
rect 327 30 385 42
rect 327 -30 339 30
rect 373 -30 385 30
rect 327 -42 385 -30
rect 505 30 563 42
rect 505 -30 517 30
rect 551 -30 563 30
rect 505 -42 563 -30
rect 683 30 741 42
rect 683 -30 695 30
rect 729 -30 741 30
rect 683 -42 741 -30
rect 861 30 919 42
rect 861 -30 873 30
rect 907 -30 919 30
rect 861 -42 919 -30
<< ndiffc >>
rect -907 -30 -873 30
rect -729 -30 -695 30
rect -551 -30 -517 30
rect -373 -30 -339 30
rect -195 -30 -161 30
rect -17 -30 17 30
rect 161 -30 195 30
rect 339 -30 373 30
rect 517 -30 551 30
rect 695 -30 729 30
rect 873 -30 907 30
<< psubdiff >>
rect -1021 182 -925 216
rect 925 182 1021 216
rect -1021 120 -987 182
rect 987 120 1021 182
rect -1021 -182 -987 -120
rect 987 -182 1021 -120
rect -1021 -216 -925 -182
rect 925 -216 1021 -182
<< psubdiffcont >>
rect -925 182 925 216
rect -1021 -120 -987 120
rect 987 -120 1021 120
rect -925 -216 925 -182
<< poly >>
rect -861 114 -741 130
rect -861 80 -845 114
rect -757 80 -741 114
rect -861 42 -741 80
rect -683 114 -563 130
rect -683 80 -667 114
rect -579 80 -563 114
rect -683 42 -563 80
rect -505 114 -385 130
rect -505 80 -489 114
rect -401 80 -385 114
rect -505 42 -385 80
rect -327 114 -207 130
rect -327 80 -311 114
rect -223 80 -207 114
rect -327 42 -207 80
rect -149 114 -29 130
rect -149 80 -133 114
rect -45 80 -29 114
rect -149 42 -29 80
rect 29 114 149 130
rect 29 80 45 114
rect 133 80 149 114
rect 29 42 149 80
rect 207 114 327 130
rect 207 80 223 114
rect 311 80 327 114
rect 207 42 327 80
rect 385 114 505 130
rect 385 80 401 114
rect 489 80 505 114
rect 385 42 505 80
rect 563 114 683 130
rect 563 80 579 114
rect 667 80 683 114
rect 563 42 683 80
rect 741 114 861 130
rect 741 80 757 114
rect 845 80 861 114
rect 741 42 861 80
rect -861 -80 -741 -42
rect -861 -114 -845 -80
rect -757 -114 -741 -80
rect -861 -130 -741 -114
rect -683 -80 -563 -42
rect -683 -114 -667 -80
rect -579 -114 -563 -80
rect -683 -130 -563 -114
rect -505 -80 -385 -42
rect -505 -114 -489 -80
rect -401 -114 -385 -80
rect -505 -130 -385 -114
rect -327 -80 -207 -42
rect -327 -114 -311 -80
rect -223 -114 -207 -80
rect -327 -130 -207 -114
rect -149 -80 -29 -42
rect -149 -114 -133 -80
rect -45 -114 -29 -80
rect -149 -130 -29 -114
rect 29 -80 149 -42
rect 29 -114 45 -80
rect 133 -114 149 -80
rect 29 -130 149 -114
rect 207 -80 327 -42
rect 207 -114 223 -80
rect 311 -114 327 -80
rect 207 -130 327 -114
rect 385 -80 505 -42
rect 385 -114 401 -80
rect 489 -114 505 -80
rect 385 -130 505 -114
rect 563 -80 683 -42
rect 563 -114 579 -80
rect 667 -114 683 -80
rect 563 -130 683 -114
rect 741 -80 861 -42
rect 741 -114 757 -80
rect 845 -114 861 -80
rect 741 -130 861 -114
<< polycont >>
rect -845 80 -757 114
rect -667 80 -579 114
rect -489 80 -401 114
rect -311 80 -223 114
rect -133 80 -45 114
rect 45 80 133 114
rect 223 80 311 114
rect 401 80 489 114
rect 579 80 667 114
rect 757 80 845 114
rect -845 -114 -757 -80
rect -667 -114 -579 -80
rect -489 -114 -401 -80
rect -311 -114 -223 -80
rect -133 -114 -45 -80
rect 45 -114 133 -80
rect 223 -114 311 -80
rect 401 -114 489 -80
rect 579 -114 667 -80
rect 757 -114 845 -80
<< locali >>
rect -1021 182 -925 216
rect 925 182 1021 216
rect -1021 120 -987 182
rect 987 120 1021 182
rect -861 80 -845 114
rect -757 80 -741 114
rect -683 80 -667 114
rect -579 80 -563 114
rect -505 80 -489 114
rect -401 80 -385 114
rect -327 80 -311 114
rect -223 80 -207 114
rect -149 80 -133 114
rect -45 80 -29 114
rect 29 80 45 114
rect 133 80 149 114
rect 207 80 223 114
rect 311 80 327 114
rect 385 80 401 114
rect 489 80 505 114
rect 563 80 579 114
rect 667 80 683 114
rect 741 80 757 114
rect 845 80 861 114
rect -907 30 -873 46
rect -907 -46 -873 -30
rect -729 30 -695 46
rect -729 -46 -695 -30
rect -551 30 -517 46
rect -551 -46 -517 -30
rect -373 30 -339 46
rect -373 -46 -339 -30
rect -195 30 -161 46
rect -195 -46 -161 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 161 30 195 46
rect 161 -46 195 -30
rect 339 30 373 46
rect 339 -46 373 -30
rect 517 30 551 46
rect 517 -46 551 -30
rect 695 30 729 46
rect 695 -46 729 -30
rect 873 30 907 46
rect 873 -46 907 -30
rect -861 -114 -845 -80
rect -757 -114 -741 -80
rect -683 -114 -667 -80
rect -579 -114 -563 -80
rect -505 -114 -489 -80
rect -401 -114 -385 -80
rect -327 -114 -311 -80
rect -223 -114 -207 -80
rect -149 -114 -133 -80
rect -45 -114 -29 -80
rect 29 -114 45 -80
rect 133 -114 149 -80
rect 207 -114 223 -80
rect 311 -114 327 -80
rect 385 -114 401 -80
rect 489 -114 505 -80
rect 563 -114 579 -80
rect 667 -114 683 -80
rect 741 -114 757 -80
rect 845 -114 861 -80
rect -1021 -182 -987 -120
rect 987 -182 1021 -120
rect -1021 -216 -925 -182
rect 925 -216 1021 -182
<< viali >>
rect -845 80 -757 114
rect -667 80 -579 114
rect -489 80 -401 114
rect -311 80 -223 114
rect -133 80 -45 114
rect 45 80 133 114
rect 223 80 311 114
rect 401 80 489 114
rect 579 80 667 114
rect 757 80 845 114
rect -907 -30 -873 30
rect -729 -30 -695 30
rect -551 -30 -517 30
rect -373 -30 -339 30
rect -195 -30 -161 30
rect -17 -30 17 30
rect 161 -30 195 30
rect 339 -30 373 30
rect 517 -30 551 30
rect 695 -30 729 30
rect 873 -30 907 30
rect -845 -114 -757 -80
rect -667 -114 -579 -80
rect -489 -114 -401 -80
rect -311 -114 -223 -80
rect -133 -114 -45 -80
rect 45 -114 133 -80
rect 223 -114 311 -80
rect 401 -114 489 -80
rect 579 -114 667 -80
rect 757 -114 845 -80
<< metal1 >>
rect -857 114 -745 120
rect -857 80 -845 114
rect -757 80 -745 114
rect -857 74 -745 80
rect -679 114 -567 120
rect -679 80 -667 114
rect -579 80 -567 114
rect -679 74 -567 80
rect -501 114 -389 120
rect -501 80 -489 114
rect -401 80 -389 114
rect -501 74 -389 80
rect -323 114 -211 120
rect -323 80 -311 114
rect -223 80 -211 114
rect -323 74 -211 80
rect -145 114 -33 120
rect -145 80 -133 114
rect -45 80 -33 114
rect -145 74 -33 80
rect 33 114 145 120
rect 33 80 45 114
rect 133 80 145 114
rect 33 74 145 80
rect 211 114 323 120
rect 211 80 223 114
rect 311 80 323 114
rect 211 74 323 80
rect 389 114 501 120
rect 389 80 401 114
rect 489 80 501 114
rect 389 74 501 80
rect 567 114 679 120
rect 567 80 579 114
rect 667 80 679 114
rect 567 74 679 80
rect 745 114 857 120
rect 745 80 757 114
rect 845 80 857 114
rect 745 74 857 80
rect -913 30 -867 42
rect -913 -30 -907 30
rect -873 -30 -867 30
rect -913 -42 -867 -30
rect -735 30 -689 42
rect -735 -30 -729 30
rect -695 -30 -689 30
rect -735 -42 -689 -30
rect -557 30 -511 42
rect -557 -30 -551 30
rect -517 -30 -511 30
rect -557 -42 -511 -30
rect -379 30 -333 42
rect -379 -30 -373 30
rect -339 -30 -333 30
rect -379 -42 -333 -30
rect -201 30 -155 42
rect -201 -30 -195 30
rect -161 -30 -155 30
rect -201 -42 -155 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 155 30 201 42
rect 155 -30 161 30
rect 195 -30 201 30
rect 155 -42 201 -30
rect 333 30 379 42
rect 333 -30 339 30
rect 373 -30 379 30
rect 333 -42 379 -30
rect 511 30 557 42
rect 511 -30 517 30
rect 551 -30 557 30
rect 511 -42 557 -30
rect 689 30 735 42
rect 689 -30 695 30
rect 729 -30 735 30
rect 689 -42 735 -30
rect 867 30 913 42
rect 867 -30 873 30
rect 907 -30 913 30
rect 867 -42 913 -30
rect -857 -80 -745 -74
rect -857 -114 -845 -80
rect -757 -114 -745 -80
rect -857 -120 -745 -114
rect -679 -80 -567 -74
rect -679 -114 -667 -80
rect -579 -114 -567 -80
rect -679 -120 -567 -114
rect -501 -80 -389 -74
rect -501 -114 -489 -80
rect -401 -114 -389 -80
rect -501 -120 -389 -114
rect -323 -80 -211 -74
rect -323 -114 -311 -80
rect -223 -114 -211 -80
rect -323 -120 -211 -114
rect -145 -80 -33 -74
rect -145 -114 -133 -80
rect -45 -114 -33 -80
rect -145 -120 -33 -114
rect 33 -80 145 -74
rect 33 -114 45 -80
rect 133 -114 145 -80
rect 33 -120 145 -114
rect 211 -80 323 -74
rect 211 -114 223 -80
rect 311 -114 323 -80
rect 211 -120 323 -114
rect 389 -80 501 -74
rect 389 -114 401 -80
rect 489 -114 501 -80
rect 389 -120 501 -114
rect 567 -80 679 -74
rect 567 -114 579 -80
rect 667 -114 679 -80
rect 567 -120 679 -114
rect 745 -80 857 -74
rect 745 -114 757 -80
rect 845 -114 857 -80
rect 745 -120 857 -114
<< properties >>
string FIXED_BBOX -1004 -199 1004 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.6 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
