** sch_path: /home/harsh/design/xschem/PLL_FOLDER/int_pfd_cp.sch
.subckt int_pfd_cp VDD cp_bias A cp_out B VSS
*.PININFO VDD:B VSS:B A:I B:I cp_bias:I cp_out:O
x1 VSS VDD A net1 net2 B pfd
x3 VDD net1 net3 VSS inverter
x2 VDD cp_bias net3 cp_out net2 VSS cp_schem
.ends

* expanding   symbol:  PLL_FOLDER/pfd.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/pfd.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/pfd.sch
.subckt pfd VSS VDD A QA QB B
*.PININFO VDD:B A:B B:B QA:B QB:B VSS:B
x1 A VDD reset VSS VSS VDD VDD QA net2 sky130_fd_sc_hd__dfrbp_2
x2 QA QB VSS VSS VDD VDD net1 sky130_fd_sc_hd__and2_2
x3 B VDD reset VSS VSS VDD VDD QB net3 sky130_fd_sc_hd__dfrbp_2
x4 net1 VSS VSS VDD VDD reset sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/harsh/design/xschem/inverter.sym
** sch_path: /home/harsh/design/xschem/inverter.sch
.subckt inverter VDD inp out VSS
*.PININFO inp:I out:O VDD:B VSS:B
x4 inp VSS VSS VDD VDD out sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  PLL_FOLDER/cp/cp_schem.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sch
.subckt cp_schem vdd cp_bias qa cp_out qb vss
*.PININFO qa:I qb:I cp_out:O vdd:B vss:B cp_bias:I
XM1 n1 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=6 nf=3 m=1
XM2 n1 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=2 nf=2 m=1
XM3 bias bias vss vss sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 m=1
XM4 n2 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=14 nf=7 m=1
XM5 n3 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.7 nf=1 m=1
XM6 cp_out qa n2 vdd sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 m=1
XM7 cp_out qb n3 vss sky130_fd_pr__nfet_01v8 L=5 W=1 nf=1 m=1
XM8 bias cp_bias vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=18 nf=9 m=1
.ends

.end
