magic
tech sky130A
magscale 1 2
timestamp 1709293017
<< error_p >>
rect -206 431 -148 437
rect -88 431 -30 437
rect 30 431 88 437
rect 148 431 206 437
rect -206 397 -194 431
rect -88 397 -76 431
rect 30 397 42 431
rect 148 397 160 431
rect -206 391 -148 397
rect -88 391 -30 397
rect 30 391 88 397
rect 148 391 206 397
rect -206 -397 -148 -391
rect -88 -397 -30 -391
rect 30 -397 88 -391
rect 148 -397 206 -391
rect -206 -431 -194 -397
rect -88 -431 -76 -397
rect 30 -431 42 -397
rect 148 -431 160 -397
rect -206 -437 -148 -431
rect -88 -437 -30 -431
rect 30 -437 88 -431
rect 148 -437 206 -431
<< nwell >>
rect -403 -569 403 569
<< pmos >>
rect -207 -350 -147 350
rect -89 -350 -29 350
rect 29 -350 89 350
rect 147 -350 207 350
<< pdiff >>
rect -265 338 -207 350
rect -265 -338 -253 338
rect -219 -338 -207 338
rect -265 -350 -207 -338
rect -147 338 -89 350
rect -147 -338 -135 338
rect -101 -338 -89 338
rect -147 -350 -89 -338
rect -29 338 29 350
rect -29 -338 -17 338
rect 17 -338 29 338
rect -29 -350 29 -338
rect 89 338 147 350
rect 89 -338 101 338
rect 135 -338 147 338
rect 89 -350 147 -338
rect 207 338 265 350
rect 207 -338 219 338
rect 253 -338 265 338
rect 207 -350 265 -338
<< pdiffc >>
rect -253 -338 -219 338
rect -135 -338 -101 338
rect -17 -338 17 338
rect 101 -338 135 338
rect 219 -338 253 338
<< nsubdiff >>
rect -367 499 -271 533
rect 271 499 367 533
rect -367 437 -333 499
rect 333 437 367 499
rect -367 -499 -333 -437
rect 333 -499 367 -437
rect -367 -533 -271 -499
rect 271 -533 367 -499
<< nsubdiffcont >>
rect -271 499 271 533
rect -367 -437 -333 437
rect 333 -437 367 437
rect -271 -533 271 -499
<< poly >>
rect -210 431 -144 447
rect -210 397 -194 431
rect -160 397 -144 431
rect -210 381 -144 397
rect -92 431 -26 447
rect -92 397 -76 431
rect -42 397 -26 431
rect -92 381 -26 397
rect 26 431 92 447
rect 26 397 42 431
rect 76 397 92 431
rect 26 381 92 397
rect 144 431 210 447
rect 144 397 160 431
rect 194 397 210 431
rect 144 381 210 397
rect -207 350 -147 381
rect -89 350 -29 381
rect 29 350 89 381
rect 147 350 207 381
rect -207 -381 -147 -350
rect -89 -381 -29 -350
rect 29 -381 89 -350
rect 147 -381 207 -350
rect -210 -397 -144 -381
rect -210 -431 -194 -397
rect -160 -431 -144 -397
rect -210 -447 -144 -431
rect -92 -397 -26 -381
rect -92 -431 -76 -397
rect -42 -431 -26 -397
rect -92 -447 -26 -431
rect 26 -397 92 -381
rect 26 -431 42 -397
rect 76 -431 92 -397
rect 26 -447 92 -431
rect 144 -397 210 -381
rect 144 -431 160 -397
rect 194 -431 210 -397
rect 144 -447 210 -431
<< polycont >>
rect -194 397 -160 431
rect -76 397 -42 431
rect 42 397 76 431
rect 160 397 194 431
rect -194 -431 -160 -397
rect -76 -431 -42 -397
rect 42 -431 76 -397
rect 160 -431 194 -397
<< locali >>
rect -367 499 -271 533
rect 271 499 367 533
rect -367 437 -333 499
rect 333 437 367 499
rect -210 397 -194 431
rect -160 397 -144 431
rect -92 397 -76 431
rect -42 397 -26 431
rect 26 397 42 431
rect 76 397 92 431
rect 144 397 160 431
rect 194 397 210 431
rect -253 338 -219 354
rect -253 -354 -219 -338
rect -135 338 -101 354
rect -135 -354 -101 -338
rect -17 338 17 354
rect -17 -354 17 -338
rect 101 338 135 354
rect 101 -354 135 -338
rect 219 338 253 354
rect 219 -354 253 -338
rect -210 -431 -194 -397
rect -160 -431 -144 -397
rect -92 -431 -76 -397
rect -42 -431 -26 -397
rect 26 -431 42 -397
rect 76 -431 92 -397
rect 144 -431 160 -397
rect 194 -431 210 -397
rect -367 -499 -333 -437
rect 333 -499 367 -437
rect -367 -533 -271 -499
rect 271 -533 367 -499
<< viali >>
rect -194 397 -160 431
rect -76 397 -42 431
rect 42 397 76 431
rect 160 397 194 431
rect -253 -338 -219 338
rect -135 -338 -101 338
rect -17 -338 17 338
rect 101 -338 135 338
rect 219 -338 253 338
rect -194 -431 -160 -397
rect -76 -431 -42 -397
rect 42 -431 76 -397
rect 160 -431 194 -397
<< metal1 >>
rect -206 431 -148 437
rect -206 397 -194 431
rect -160 397 -148 431
rect -206 391 -148 397
rect -88 431 -30 437
rect -88 397 -76 431
rect -42 397 -30 431
rect -88 391 -30 397
rect 30 431 88 437
rect 30 397 42 431
rect 76 397 88 431
rect 30 391 88 397
rect 148 431 206 437
rect 148 397 160 431
rect 194 397 206 431
rect 148 391 206 397
rect -259 338 -213 350
rect -259 -338 -253 338
rect -219 -338 -213 338
rect -259 -350 -213 -338
rect -141 338 -95 350
rect -141 -338 -135 338
rect -101 -338 -95 338
rect -141 -350 -95 -338
rect -23 338 23 350
rect -23 -338 -17 338
rect 17 -338 23 338
rect -23 -350 23 -338
rect 95 338 141 350
rect 95 -338 101 338
rect 135 -338 141 338
rect 95 -350 141 -338
rect 213 338 259 350
rect 213 -338 219 338
rect 253 -338 259 338
rect 213 -350 259 -338
rect -206 -397 -148 -391
rect -206 -431 -194 -397
rect -160 -431 -148 -397
rect -206 -437 -148 -431
rect -88 -397 -30 -391
rect -88 -431 -76 -397
rect -42 -431 -30 -397
rect -88 -437 -30 -431
rect 30 -397 88 -391
rect 30 -431 42 -397
rect 76 -431 88 -397
rect 30 -437 88 -431
rect 148 -397 206 -391
rect 148 -431 160 -397
rect 194 -431 206 -397
rect 148 -437 206 -431
<< properties >>
string FIXED_BBOX -350 -516 350 516
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.5 l 0.3 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
