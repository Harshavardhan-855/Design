magic
tech sky130A
timestamp 1708417395
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
use sky130_fd_sc_hd__inv_4  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform 1 0 631 0 1 101
box -19 -24 249 296
use sky130_fd_sc_hd__inv_4  x4
timestamp 1705271942
transform 1 0 -430 0 1 152
box -19 -24 249 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 inp
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 out
port 3 nsew
<< end >>
