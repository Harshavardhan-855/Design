magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< error_p >>
rect -560 114 -502 120
rect -442 114 -384 120
rect -324 114 -266 120
rect -206 114 -148 120
rect -88 114 -30 120
rect 30 114 88 120
rect 148 114 206 120
rect 266 114 324 120
rect 384 114 442 120
rect 502 114 560 120
rect -560 80 -548 114
rect -442 80 -430 114
rect -324 80 -312 114
rect -206 80 -194 114
rect -88 80 -76 114
rect 30 80 42 114
rect 148 80 160 114
rect 266 80 278 114
rect 384 80 396 114
rect 502 80 514 114
rect -560 74 -502 80
rect -442 74 -384 80
rect -324 74 -266 80
rect -206 74 -148 80
rect -88 74 -30 80
rect 30 74 88 80
rect 148 74 206 80
rect 266 74 324 80
rect 384 74 442 80
rect 502 74 560 80
rect -560 -80 -502 -74
rect -442 -80 -384 -74
rect -324 -80 -266 -74
rect -206 -80 -148 -74
rect -88 -80 -30 -74
rect 30 -80 88 -74
rect 148 -80 206 -74
rect 266 -80 324 -74
rect 384 -80 442 -74
rect 502 -80 560 -74
rect -560 -114 -548 -80
rect -442 -114 -430 -80
rect -324 -114 -312 -80
rect -206 -114 -194 -80
rect -88 -114 -76 -80
rect 30 -114 42 -80
rect 148 -114 160 -80
rect 266 -114 278 -80
rect 384 -114 396 -80
rect 502 -114 514 -80
rect -560 -120 -502 -114
rect -442 -120 -384 -114
rect -324 -120 -266 -114
rect -206 -120 -148 -114
rect -88 -120 -30 -114
rect 30 -120 88 -114
rect 148 -120 206 -114
rect 266 -120 324 -114
rect 384 -120 442 -114
rect 502 -120 560 -114
<< pwell >>
rect -757 -252 757 252
<< nmos >>
rect -561 -42 -501 42
rect -443 -42 -383 42
rect -325 -42 -265 42
rect -207 -42 -147 42
rect -89 -42 -29 42
rect 29 -42 89 42
rect 147 -42 207 42
rect 265 -42 325 42
rect 383 -42 443 42
rect 501 -42 561 42
<< ndiff >>
rect -619 30 -561 42
rect -619 -30 -607 30
rect -573 -30 -561 30
rect -619 -42 -561 -30
rect -501 30 -443 42
rect -501 -30 -489 30
rect -455 -30 -443 30
rect -501 -42 -443 -30
rect -383 30 -325 42
rect -383 -30 -371 30
rect -337 -30 -325 30
rect -383 -42 -325 -30
rect -265 30 -207 42
rect -265 -30 -253 30
rect -219 -30 -207 30
rect -265 -42 -207 -30
rect -147 30 -89 42
rect -147 -30 -135 30
rect -101 -30 -89 30
rect -147 -42 -89 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 89 30 147 42
rect 89 -30 101 30
rect 135 -30 147 30
rect 89 -42 147 -30
rect 207 30 265 42
rect 207 -30 219 30
rect 253 -30 265 30
rect 207 -42 265 -30
rect 325 30 383 42
rect 325 -30 337 30
rect 371 -30 383 30
rect 325 -42 383 -30
rect 443 30 501 42
rect 443 -30 455 30
rect 489 -30 501 30
rect 443 -42 501 -30
rect 561 30 619 42
rect 561 -30 573 30
rect 607 -30 619 30
rect 561 -42 619 -30
<< ndiffc >>
rect -607 -30 -573 30
rect -489 -30 -455 30
rect -371 -30 -337 30
rect -253 -30 -219 30
rect -135 -30 -101 30
rect -17 -30 17 30
rect 101 -30 135 30
rect 219 -30 253 30
rect 337 -30 371 30
rect 455 -30 489 30
rect 573 -30 607 30
<< psubdiff >>
rect -721 182 -625 216
rect 625 182 721 216
rect -721 120 -687 182
rect 687 120 721 182
rect -721 -182 -687 -120
rect 687 -182 721 -120
rect -721 -216 -625 -182
rect 625 -216 721 -182
<< psubdiffcont >>
rect -625 182 625 216
rect -721 -120 -687 120
rect 687 -120 721 120
rect -625 -216 625 -182
<< poly >>
rect -564 114 -498 130
rect -564 80 -548 114
rect -514 80 -498 114
rect -564 64 -498 80
rect -446 114 -380 130
rect -446 80 -430 114
rect -396 80 -380 114
rect -446 64 -380 80
rect -328 114 -262 130
rect -328 80 -312 114
rect -278 80 -262 114
rect -328 64 -262 80
rect -210 114 -144 130
rect -210 80 -194 114
rect -160 80 -144 114
rect -210 64 -144 80
rect -92 114 -26 130
rect -92 80 -76 114
rect -42 80 -26 114
rect -92 64 -26 80
rect 26 114 92 130
rect 26 80 42 114
rect 76 80 92 114
rect 26 64 92 80
rect 144 114 210 130
rect 144 80 160 114
rect 194 80 210 114
rect 144 64 210 80
rect 262 114 328 130
rect 262 80 278 114
rect 312 80 328 114
rect 262 64 328 80
rect 380 114 446 130
rect 380 80 396 114
rect 430 80 446 114
rect 380 64 446 80
rect 498 114 564 130
rect 498 80 514 114
rect 548 80 564 114
rect 498 64 564 80
rect -561 42 -501 64
rect -443 42 -383 64
rect -325 42 -265 64
rect -207 42 -147 64
rect -89 42 -29 64
rect 29 42 89 64
rect 147 42 207 64
rect 265 42 325 64
rect 383 42 443 64
rect 501 42 561 64
rect -561 -64 -501 -42
rect -443 -64 -383 -42
rect -325 -64 -265 -42
rect -207 -64 -147 -42
rect -89 -64 -29 -42
rect 29 -64 89 -42
rect 147 -64 207 -42
rect 265 -64 325 -42
rect 383 -64 443 -42
rect 501 -64 561 -42
rect -564 -80 -498 -64
rect -564 -114 -548 -80
rect -514 -114 -498 -80
rect -564 -130 -498 -114
rect -446 -80 -380 -64
rect -446 -114 -430 -80
rect -396 -114 -380 -80
rect -446 -130 -380 -114
rect -328 -80 -262 -64
rect -328 -114 -312 -80
rect -278 -114 -262 -80
rect -328 -130 -262 -114
rect -210 -80 -144 -64
rect -210 -114 -194 -80
rect -160 -114 -144 -80
rect -210 -130 -144 -114
rect -92 -80 -26 -64
rect -92 -114 -76 -80
rect -42 -114 -26 -80
rect -92 -130 -26 -114
rect 26 -80 92 -64
rect 26 -114 42 -80
rect 76 -114 92 -80
rect 26 -130 92 -114
rect 144 -80 210 -64
rect 144 -114 160 -80
rect 194 -114 210 -80
rect 144 -130 210 -114
rect 262 -80 328 -64
rect 262 -114 278 -80
rect 312 -114 328 -80
rect 262 -130 328 -114
rect 380 -80 446 -64
rect 380 -114 396 -80
rect 430 -114 446 -80
rect 380 -130 446 -114
rect 498 -80 564 -64
rect 498 -114 514 -80
rect 548 -114 564 -80
rect 498 -130 564 -114
<< polycont >>
rect -548 80 -514 114
rect -430 80 -396 114
rect -312 80 -278 114
rect -194 80 -160 114
rect -76 80 -42 114
rect 42 80 76 114
rect 160 80 194 114
rect 278 80 312 114
rect 396 80 430 114
rect 514 80 548 114
rect -548 -114 -514 -80
rect -430 -114 -396 -80
rect -312 -114 -278 -80
rect -194 -114 -160 -80
rect -76 -114 -42 -80
rect 42 -114 76 -80
rect 160 -114 194 -80
rect 278 -114 312 -80
rect 396 -114 430 -80
rect 514 -114 548 -80
<< locali >>
rect -721 182 -625 216
rect 625 182 721 216
rect -721 120 -687 182
rect 687 120 721 182
rect -564 80 -548 114
rect -514 80 -498 114
rect -446 80 -430 114
rect -396 80 -380 114
rect -328 80 -312 114
rect -278 80 -262 114
rect -210 80 -194 114
rect -160 80 -144 114
rect -92 80 -76 114
rect -42 80 -26 114
rect 26 80 42 114
rect 76 80 92 114
rect 144 80 160 114
rect 194 80 210 114
rect 262 80 278 114
rect 312 80 328 114
rect 380 80 396 114
rect 430 80 446 114
rect 498 80 514 114
rect 548 80 564 114
rect -607 30 -573 46
rect -607 -46 -573 -30
rect -489 30 -455 46
rect -489 -46 -455 -30
rect -371 30 -337 46
rect -371 -46 -337 -30
rect -253 30 -219 46
rect -253 -46 -219 -30
rect -135 30 -101 46
rect -135 -46 -101 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 101 30 135 46
rect 101 -46 135 -30
rect 219 30 253 46
rect 219 -46 253 -30
rect 337 30 371 46
rect 337 -46 371 -30
rect 455 30 489 46
rect 455 -46 489 -30
rect 573 30 607 46
rect 573 -46 607 -30
rect -564 -114 -548 -80
rect -514 -114 -498 -80
rect -446 -114 -430 -80
rect -396 -114 -380 -80
rect -328 -114 -312 -80
rect -278 -114 -262 -80
rect -210 -114 -194 -80
rect -160 -114 -144 -80
rect -92 -114 -76 -80
rect -42 -114 -26 -80
rect 26 -114 42 -80
rect 76 -114 92 -80
rect 144 -114 160 -80
rect 194 -114 210 -80
rect 262 -114 278 -80
rect 312 -114 328 -80
rect 380 -114 396 -80
rect 430 -114 446 -80
rect 498 -114 514 -80
rect 548 -114 564 -80
rect -721 -182 -687 -120
rect 687 -182 721 -120
rect -721 -216 -625 -182
rect 625 -216 721 -182
<< viali >>
rect -548 80 -514 114
rect -430 80 -396 114
rect -312 80 -278 114
rect -194 80 -160 114
rect -76 80 -42 114
rect 42 80 76 114
rect 160 80 194 114
rect 278 80 312 114
rect 396 80 430 114
rect 514 80 548 114
rect -607 -30 -573 30
rect -489 -30 -455 30
rect -371 -30 -337 30
rect -253 -30 -219 30
rect -135 -30 -101 30
rect -17 -30 17 30
rect 101 -30 135 30
rect 219 -30 253 30
rect 337 -30 371 30
rect 455 -30 489 30
rect 573 -30 607 30
rect -548 -114 -514 -80
rect -430 -114 -396 -80
rect -312 -114 -278 -80
rect -194 -114 -160 -80
rect -76 -114 -42 -80
rect 42 -114 76 -80
rect 160 -114 194 -80
rect 278 -114 312 -80
rect 396 -114 430 -80
rect 514 -114 548 -80
<< metal1 >>
rect -560 114 -502 120
rect -560 80 -548 114
rect -514 80 -502 114
rect -560 74 -502 80
rect -442 114 -384 120
rect -442 80 -430 114
rect -396 80 -384 114
rect -442 74 -384 80
rect -324 114 -266 120
rect -324 80 -312 114
rect -278 80 -266 114
rect -324 74 -266 80
rect -206 114 -148 120
rect -206 80 -194 114
rect -160 80 -148 114
rect -206 74 -148 80
rect -88 114 -30 120
rect -88 80 -76 114
rect -42 80 -30 114
rect -88 74 -30 80
rect 30 114 88 120
rect 30 80 42 114
rect 76 80 88 114
rect 30 74 88 80
rect 148 114 206 120
rect 148 80 160 114
rect 194 80 206 114
rect 148 74 206 80
rect 266 114 324 120
rect 266 80 278 114
rect 312 80 324 114
rect 266 74 324 80
rect 384 114 442 120
rect 384 80 396 114
rect 430 80 442 114
rect 384 74 442 80
rect 502 114 560 120
rect 502 80 514 114
rect 548 80 560 114
rect 502 74 560 80
rect -613 30 -567 42
rect -613 -30 -607 30
rect -573 -30 -567 30
rect -613 -42 -567 -30
rect -495 30 -449 42
rect -495 -30 -489 30
rect -455 -30 -449 30
rect -495 -42 -449 -30
rect -377 30 -331 42
rect -377 -30 -371 30
rect -337 -30 -331 30
rect -377 -42 -331 -30
rect -259 30 -213 42
rect -259 -30 -253 30
rect -219 -30 -213 30
rect -259 -42 -213 -30
rect -141 30 -95 42
rect -141 -30 -135 30
rect -101 -30 -95 30
rect -141 -42 -95 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 95 30 141 42
rect 95 -30 101 30
rect 135 -30 141 30
rect 95 -42 141 -30
rect 213 30 259 42
rect 213 -30 219 30
rect 253 -30 259 30
rect 213 -42 259 -30
rect 331 30 377 42
rect 331 -30 337 30
rect 371 -30 377 30
rect 331 -42 377 -30
rect 449 30 495 42
rect 449 -30 455 30
rect 489 -30 495 30
rect 449 -42 495 -30
rect 567 30 613 42
rect 567 -30 573 30
rect 607 -30 613 30
rect 567 -42 613 -30
rect -560 -80 -502 -74
rect -560 -114 -548 -80
rect -514 -114 -502 -80
rect -560 -120 -502 -114
rect -442 -80 -384 -74
rect -442 -114 -430 -80
rect -396 -114 -384 -80
rect -442 -120 -384 -114
rect -324 -80 -266 -74
rect -324 -114 -312 -80
rect -278 -114 -266 -80
rect -324 -120 -266 -114
rect -206 -80 -148 -74
rect -206 -114 -194 -80
rect -160 -114 -148 -80
rect -206 -120 -148 -114
rect -88 -80 -30 -74
rect -88 -114 -76 -80
rect -42 -114 -30 -80
rect -88 -120 -30 -114
rect 30 -80 88 -74
rect 30 -114 42 -80
rect 76 -114 88 -80
rect 30 -120 88 -114
rect 148 -80 206 -74
rect 148 -114 160 -80
rect 194 -114 206 -80
rect 148 -120 206 -114
rect 266 -80 324 -74
rect 266 -114 278 -80
rect 312 -114 324 -80
rect 266 -120 324 -114
rect 384 -80 442 -74
rect 384 -114 396 -80
rect 430 -114 442 -80
rect 384 -120 442 -114
rect 502 -80 560 -74
rect 502 -114 514 -80
rect 548 -114 560 -80
rect 502 -120 560 -114
<< properties >>
string FIXED_BBOX -704 -199 704 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
