** UNTITLED-9 flat netlist

*--------BEGIN_X1->INT_PFD_CP
*.PININFO VDD:B VSS:B A:I B:I CP_BIAS:I CP_OUT:O
*--------BEGIN_X1_X1->PFD
*.PININFO VDD:B A:B B:B QA:B QB:B VSS:B
*--------BEGIN_X1_X1_X1->SKY130_FD_SC_HD__DFRBP_2
X1_X1_X1 NET3 NET1 X1_X1_RESET X1_NET4 X1_NET4 NET1 NET1 X1_NET1 X1_X1_NET2  SKY130_FD_SC_HD__DFRBP_2
*--------END___X1_X1_X1->SKY130_FD_SC_HD__DFRBP_2
*--------BEGIN_X1_X1_X2->SKY130_FD_SC_HD__AND2_2
X2_X1_X1 X1_NET1 X1_NET3 X1_NET4 X1_NET4 NET1 NET1 X1_X1_NET1  SKY130_FD_SC_HD__AND2_2
*--------END___X1_X1_X2->SKY130_FD_SC_HD__AND2_2
*--------BEGIN_X1_X1_X3->SKY130_FD_SC_HD__DFRBP_2
X3_X1_X1 NET5 NET1 X1_X1_RESET X1_NET4 X1_NET4 NET1 NET1 X1_NET3 X1_X1_NET3  SKY130_FD_SC_HD__DFRBP_2
*--------END___X1_X1_X3->SKY130_FD_SC_HD__DFRBP_2
*--------BEGIN_X1_X1_X4->SKY130_FD_SC_HD__INV_4
X4_X1_X1 X1_X1_NET1 X1_NET4 X1_NET4 NET1 NET1 X1_X1_RESET  SKY130_FD_SC_HD__INV_4
*--------END___X1_X1_X4->SKY130_FD_SC_HD__INV_4
*--------END___X1_X1->PFD
*--------BEGIN_X1_X2->CP_SCHEM

*--------END___X1_X2->CP_SCHEM
*--------BEGIN_X1_X3->INVERTER
*.PININFO INP:I OUT:O VDD:B VSS:B
*--------BEGIN_X1_X3_X4->SKY130_FD_SC_HD__INV_4
X4_X1_X3 X1_NET1 NET6 NET6 NET1 NET1 X1_NET2  SKY130_FD_SC_HD__INV_4
*--------END___X1_X3_X4->SKY130_FD_SC_HD__INV_4
*--------END___X1_X3->INVERTER
*  X1 -       IS MISSING !!!!
*--------END___X1->INT_PFD_CP
.end
