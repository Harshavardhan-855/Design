** sch_path: /home/harsh/design/xschem/PLL_FOLDER/top_pll.sch
.subckt top_pll Ref_sig i_bias vco_out vdd vss
*.PININFO Ref_sig:I i_bias:I vco_out:O vdd:B vss:B
x1 vss vdd Ref_sig net1 net2 net4 pfd
x3 vdd vco_out net3 vss vco
x4 vdd net1 net5 vss inverter
x5 vdd net6 net4 net7 vco_out vss divider_3N
x2 vdd i_bias net5 net3 net2 vss cp_schem
.ends

* expanding   symbol:  PLL_FOLDER/pfd.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/pfd.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/pfd.sch
.subckt pfd VSS VDD A QA QB B
*.PININFO VDD:B A:B B:B QA:B QB:B VSS:B
x1 A VDD reset VSS VSS VDD VDD QA net2 sky130_fd_sc_hd__dfrbp_2
x2 QA QB VSS VSS VDD VDD net1 sky130_fd_sc_hd__and2_2
x3 B VDD reset VSS VSS VDD VDD QB net3 sky130_fd_sc_hd__dfrbp_2
x4 net1 VSS VSS VDD VDD reset sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  PLL_FOLDER/vco/vco.sym # of pins=4
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/vco/vco.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/vco/vco.sch
.subckt vco vdd out vctrl vss
*.PININFO vdd:B vss:B out:B vctrl:B
XM1 net1 vctrl vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=30 nf=5 m=1
XM2 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=90 nf=5 m=1
XM3 net4 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=80 nf=10 m=1
XM4 net3 out net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=80 nf=10 m=1
XM5 net2 vctrl vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=30 nf=10 m=1
XM6 net3 out net2 vss sky130_fd_pr__nfet_01v8 L=0.15 W=30 nf=10 m=1
XM7 net7 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=160 nf=20 m=1
XM8 net6 net3 net7 net7 sky130_fd_pr__pfet_01v8 L=0.15 W=160 nf=20 m=1
XM9 net5 vctrl vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=60 nf=20 m=1
XM10 net6 net3 net5 vss sky130_fd_pr__nfet_01v8 L=0.15 W=60 nf=20 m=1
XM11 net9 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=240 nf=30 m=1
XM12 out net6 net9 net9 sky130_fd_pr__pfet_01v8 L=0.15 W=240 nf=30 m=1
XM13 net8 vctrl vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=90 nf=30 m=1
XM14 out net6 net8 vss sky130_fd_pr__nfet_01v8 L=0.15 W=90 nf=30 m=1
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/harsh/design/xschem/inverter.sym
** sch_path: /home/harsh/design/xschem/inverter.sch
.subckt inverter VDD inp out VSS
*.PININFO inp:I out:O VDD:B VSS:B
x4 inp VSS VSS VDD VDD out sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  PLL_FOLDER/divider/divider_3N.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/divider/divider_3N.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/divider/divider_3N.sch
.subckt divider_3N vdd out_b out_c out_a clock vss
*.PININFO clock:I out_a:O out_b:O out_c:O vdd:B vss:B
x3 clock net1 VSS VSS VDD VDD out_a net1 sky130_fd_sc_hd__dfxbp_2
x1 net1 net2 VSS VSS VDD VDD out_b net2 sky130_fd_sc_hd__dfxbp_2
x2 net2 net3 VSS VSS VDD VDD out_c net3 sky130_fd_sc_hd__dfxbp_2
.ends


* expanding   symbol:  PLL_FOLDER/cp/cp_schem.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sch
.subckt cp_schem vdd cp_bias qa cp_out qb vss
*.PININFO qa:I qb:I cp_out:O vdd:B vss:B cp_bias:I
XM1 n1 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=6 nf=3 m=1
XM2 n1 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=2 nf=2 m=1
XM3 bias bias vss vss sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 m=1
XM4 n2 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=14 nf=7 m=1
XM5 n3 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.7 nf=1 m=1
XM6 cp_out qa n2 vdd sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 m=1
XM7 cp_out qb n3 vss sky130_fd_pr__nfet_01v8 L=5 W=1 nf=1 m=1
XM8 bias cp_bias vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=18 nf=9 m=1
.ends

.end
