magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -365 161 -307 167
rect -173 161 -115 167
rect 19 161 77 167
rect 211 161 269 167
rect 403 161 461 167
rect -365 127 -353 161
rect -173 127 -161 161
rect 19 127 31 161
rect 211 127 223 161
rect 403 127 415 161
rect -365 121 -307 127
rect -173 121 -115 127
rect 19 121 77 127
rect 211 121 269 127
rect 403 121 461 127
rect -461 -127 -403 -121
rect -269 -127 -211 -121
rect -77 -127 -19 -121
rect 115 -127 173 -121
rect 307 -127 365 -121
rect -461 -161 -449 -127
rect -269 -161 -257 -127
rect -77 -161 -65 -127
rect 115 -161 127 -127
rect 307 -161 319 -127
rect -461 -167 -403 -161
rect -269 -167 -211 -161
rect -77 -167 -19 -161
rect 115 -167 173 -161
rect 307 -167 365 -161
<< nwell >>
rect -647 -299 647 299
<< pmos >>
rect -447 -80 -417 80
rect -351 -80 -321 80
rect -255 -80 -225 80
rect -159 -80 -129 80
rect -63 -80 -33 80
rect 33 -80 63 80
rect 129 -80 159 80
rect 225 -80 255 80
rect 321 -80 351 80
rect 417 -80 447 80
<< pdiff >>
rect -509 68 -447 80
rect -509 -68 -497 68
rect -463 -68 -447 68
rect -509 -80 -447 -68
rect -417 68 -351 80
rect -417 -68 -401 68
rect -367 -68 -351 68
rect -417 -80 -351 -68
rect -321 68 -255 80
rect -321 -68 -305 68
rect -271 -68 -255 68
rect -321 -80 -255 -68
rect -225 68 -159 80
rect -225 -68 -209 68
rect -175 -68 -159 68
rect -225 -80 -159 -68
rect -129 68 -63 80
rect -129 -68 -113 68
rect -79 -68 -63 68
rect -129 -80 -63 -68
rect -33 68 33 80
rect -33 -68 -17 68
rect 17 -68 33 68
rect -33 -80 33 -68
rect 63 68 129 80
rect 63 -68 79 68
rect 113 -68 129 68
rect 63 -80 129 -68
rect 159 68 225 80
rect 159 -68 175 68
rect 209 -68 225 68
rect 159 -80 225 -68
rect 255 68 321 80
rect 255 -68 271 68
rect 305 -68 321 68
rect 255 -80 321 -68
rect 351 68 417 80
rect 351 -68 367 68
rect 401 -68 417 68
rect 351 -80 417 -68
rect 447 68 509 80
rect 447 -68 463 68
rect 497 -68 509 68
rect 447 -80 509 -68
<< pdiffc >>
rect -497 -68 -463 68
rect -401 -68 -367 68
rect -305 -68 -271 68
rect -209 -68 -175 68
rect -113 -68 -79 68
rect -17 -68 17 68
rect 79 -68 113 68
rect 175 -68 209 68
rect 271 -68 305 68
rect 367 -68 401 68
rect 463 -68 497 68
<< nsubdiff >>
rect -611 229 -515 263
rect 515 229 611 263
rect -611 167 -577 229
rect 577 167 611 229
rect -611 -229 -577 -167
rect 577 -229 611 -167
rect -611 -263 -515 -229
rect 515 -263 611 -229
<< nsubdiffcont >>
rect -515 229 515 263
rect -611 -167 -577 167
rect 577 -167 611 167
rect -515 -263 515 -229
<< poly >>
rect -369 161 -303 177
rect -369 127 -353 161
rect -319 127 -303 161
rect -369 111 -303 127
rect -177 161 -111 177
rect -177 127 -161 161
rect -127 127 -111 161
rect -177 111 -111 127
rect 15 161 81 177
rect 15 127 31 161
rect 65 127 81 161
rect 15 111 81 127
rect 207 161 273 177
rect 207 127 223 161
rect 257 127 273 161
rect 207 111 273 127
rect 399 161 465 177
rect 399 127 415 161
rect 449 127 465 161
rect 399 111 465 127
rect -447 80 -417 106
rect -351 80 -321 111
rect -255 80 -225 106
rect -159 80 -129 111
rect -63 80 -33 106
rect 33 80 63 111
rect 129 80 159 106
rect 225 80 255 111
rect 321 80 351 106
rect 417 80 447 111
rect -447 -111 -417 -80
rect -351 -106 -321 -80
rect -255 -111 -225 -80
rect -159 -106 -129 -80
rect -63 -111 -33 -80
rect 33 -106 63 -80
rect 129 -111 159 -80
rect 225 -106 255 -80
rect 321 -111 351 -80
rect 417 -106 447 -80
rect -465 -127 -399 -111
rect -465 -161 -449 -127
rect -415 -161 -399 -127
rect -465 -177 -399 -161
rect -273 -127 -207 -111
rect -273 -161 -257 -127
rect -223 -161 -207 -127
rect -273 -177 -207 -161
rect -81 -127 -15 -111
rect -81 -161 -65 -127
rect -31 -161 -15 -127
rect -81 -177 -15 -161
rect 111 -127 177 -111
rect 111 -161 127 -127
rect 161 -161 177 -127
rect 111 -177 177 -161
rect 303 -127 369 -111
rect 303 -161 319 -127
rect 353 -161 369 -127
rect 303 -177 369 -161
<< polycont >>
rect -353 127 -319 161
rect -161 127 -127 161
rect 31 127 65 161
rect 223 127 257 161
rect 415 127 449 161
rect -449 -161 -415 -127
rect -257 -161 -223 -127
rect -65 -161 -31 -127
rect 127 -161 161 -127
rect 319 -161 353 -127
<< locali >>
rect -611 229 -515 263
rect 515 229 611 263
rect -611 167 -577 229
rect 577 167 611 229
rect -369 127 -353 161
rect -319 127 -303 161
rect -177 127 -161 161
rect -127 127 -111 161
rect 15 127 31 161
rect 65 127 81 161
rect 207 127 223 161
rect 257 127 273 161
rect 399 127 415 161
rect 449 127 465 161
rect -497 68 -463 84
rect -497 -84 -463 -68
rect -401 68 -367 84
rect -401 -84 -367 -68
rect -305 68 -271 84
rect -305 -84 -271 -68
rect -209 68 -175 84
rect -209 -84 -175 -68
rect -113 68 -79 84
rect -113 -84 -79 -68
rect -17 68 17 84
rect -17 -84 17 -68
rect 79 68 113 84
rect 79 -84 113 -68
rect 175 68 209 84
rect 175 -84 209 -68
rect 271 68 305 84
rect 271 -84 305 -68
rect 367 68 401 84
rect 367 -84 401 -68
rect 463 68 497 84
rect 463 -84 497 -68
rect -465 -161 -449 -127
rect -415 -161 -399 -127
rect -273 -161 -257 -127
rect -223 -161 -207 -127
rect -81 -161 -65 -127
rect -31 -161 -15 -127
rect 111 -161 127 -127
rect 161 -161 177 -127
rect 303 -161 319 -127
rect 353 -161 369 -127
rect -611 -229 -577 -167
rect 577 -229 611 -167
rect -611 -263 -515 -229
rect 515 -263 611 -229
<< viali >>
rect -353 127 -319 161
rect -161 127 -127 161
rect 31 127 65 161
rect 223 127 257 161
rect 415 127 449 161
rect -497 -68 -463 68
rect -401 -68 -367 68
rect -305 -68 -271 68
rect -209 -68 -175 68
rect -113 -68 -79 68
rect -17 -68 17 68
rect 79 -68 113 68
rect 175 -68 209 68
rect 271 -68 305 68
rect 367 -68 401 68
rect 463 -68 497 68
rect -449 -161 -415 -127
rect -257 -161 -223 -127
rect -65 -161 -31 -127
rect 127 -161 161 -127
rect 319 -161 353 -127
<< metal1 >>
rect -365 161 -307 167
rect -365 127 -353 161
rect -319 127 -307 161
rect -365 121 -307 127
rect -173 161 -115 167
rect -173 127 -161 161
rect -127 127 -115 161
rect -173 121 -115 127
rect 19 161 77 167
rect 19 127 31 161
rect 65 127 77 161
rect 19 121 77 127
rect 211 161 269 167
rect 211 127 223 161
rect 257 127 269 161
rect 211 121 269 127
rect 403 161 461 167
rect 403 127 415 161
rect 449 127 461 161
rect 403 121 461 127
rect -503 68 -457 80
rect -503 -68 -497 68
rect -463 -68 -457 68
rect -503 -80 -457 -68
rect -407 68 -361 80
rect -407 -68 -401 68
rect -367 -68 -361 68
rect -407 -80 -361 -68
rect -311 68 -265 80
rect -311 -68 -305 68
rect -271 -68 -265 68
rect -311 -80 -265 -68
rect -215 68 -169 80
rect -215 -68 -209 68
rect -175 -68 -169 68
rect -215 -80 -169 -68
rect -119 68 -73 80
rect -119 -68 -113 68
rect -79 -68 -73 68
rect -119 -80 -73 -68
rect -23 68 23 80
rect -23 -68 -17 68
rect 17 -68 23 68
rect -23 -80 23 -68
rect 73 68 119 80
rect 73 -68 79 68
rect 113 -68 119 68
rect 73 -80 119 -68
rect 169 68 215 80
rect 169 -68 175 68
rect 209 -68 215 68
rect 169 -80 215 -68
rect 265 68 311 80
rect 265 -68 271 68
rect 305 -68 311 68
rect 265 -80 311 -68
rect 361 68 407 80
rect 361 -68 367 68
rect 401 -68 407 68
rect 361 -80 407 -68
rect 457 68 503 80
rect 457 -68 463 68
rect 497 -68 503 68
rect 457 -80 503 -68
rect -461 -127 -403 -121
rect -461 -161 -449 -127
rect -415 -161 -403 -127
rect -461 -167 -403 -161
rect -269 -127 -211 -121
rect -269 -161 -257 -127
rect -223 -161 -211 -127
rect -269 -167 -211 -161
rect -77 -127 -19 -121
rect -77 -161 -65 -127
rect -31 -161 -19 -127
rect -77 -167 -19 -161
rect 115 -127 173 -121
rect 115 -161 127 -127
rect 161 -161 173 -127
rect 115 -167 173 -161
rect 307 -127 365 -121
rect 307 -161 319 -127
rect 353 -161 365 -127
rect 307 -167 365 -161
<< properties >>
string FIXED_BBOX -594 -246 594 246
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
