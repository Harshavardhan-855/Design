magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< error_p >>
rect -855 1272 -797 1278
rect -737 1272 -679 1278
rect -619 1272 -561 1278
rect -501 1272 -443 1278
rect -383 1272 -325 1278
rect -265 1272 -207 1278
rect -147 1272 -89 1278
rect -29 1272 29 1278
rect 89 1272 147 1278
rect 207 1272 265 1278
rect 325 1272 383 1278
rect 443 1272 501 1278
rect 561 1272 619 1278
rect 679 1272 737 1278
rect 797 1272 855 1278
rect -855 1238 -843 1272
rect -737 1238 -725 1272
rect -619 1238 -607 1272
rect -501 1238 -489 1272
rect -383 1238 -371 1272
rect -265 1238 -253 1272
rect -147 1238 -135 1272
rect -29 1238 -17 1272
rect 89 1238 101 1272
rect 207 1238 219 1272
rect 325 1238 337 1272
rect 443 1238 455 1272
rect 561 1238 573 1272
rect 679 1238 691 1272
rect 797 1238 809 1272
rect -855 1232 -797 1238
rect -737 1232 -679 1238
rect -619 1232 -561 1238
rect -501 1232 -443 1238
rect -383 1232 -325 1238
rect -265 1232 -207 1238
rect -147 1232 -89 1238
rect -29 1232 29 1238
rect 89 1232 147 1238
rect 207 1232 265 1238
rect 325 1232 383 1238
rect 443 1232 501 1238
rect 561 1232 619 1238
rect 679 1232 737 1238
rect 797 1232 855 1238
rect -855 -1238 -797 -1232
rect -737 -1238 -679 -1232
rect -619 -1238 -561 -1232
rect -501 -1238 -443 -1232
rect -383 -1238 -325 -1232
rect -265 -1238 -207 -1232
rect -147 -1238 -89 -1232
rect -29 -1238 29 -1232
rect 89 -1238 147 -1232
rect 207 -1238 265 -1232
rect 325 -1238 383 -1232
rect 443 -1238 501 -1232
rect 561 -1238 619 -1232
rect 679 -1238 737 -1232
rect 797 -1238 855 -1232
rect -855 -1272 -843 -1238
rect -737 -1272 -725 -1238
rect -619 -1272 -607 -1238
rect -501 -1272 -489 -1238
rect -383 -1272 -371 -1238
rect -265 -1272 -253 -1238
rect -147 -1272 -135 -1238
rect -29 -1272 -17 -1238
rect 89 -1272 101 -1238
rect 207 -1272 219 -1238
rect 325 -1272 337 -1238
rect 443 -1272 455 -1238
rect 561 -1272 573 -1238
rect 679 -1272 691 -1238
rect 797 -1272 809 -1238
rect -855 -1278 -797 -1272
rect -737 -1278 -679 -1272
rect -619 -1278 -561 -1272
rect -501 -1278 -443 -1272
rect -383 -1278 -325 -1272
rect -265 -1278 -207 -1272
rect -147 -1278 -89 -1272
rect -29 -1278 29 -1272
rect 89 -1278 147 -1272
rect 207 -1278 265 -1272
rect 325 -1278 383 -1272
rect 443 -1278 501 -1272
rect 561 -1278 619 -1272
rect 679 -1278 737 -1272
rect 797 -1278 855 -1272
<< pwell >>
rect -1052 -1410 1052 1410
<< nmos >>
rect -856 -1200 -796 1200
rect -738 -1200 -678 1200
rect -620 -1200 -560 1200
rect -502 -1200 -442 1200
rect -384 -1200 -324 1200
rect -266 -1200 -206 1200
rect -148 -1200 -88 1200
rect -30 -1200 30 1200
rect 88 -1200 148 1200
rect 206 -1200 266 1200
rect 324 -1200 384 1200
rect 442 -1200 502 1200
rect 560 -1200 620 1200
rect 678 -1200 738 1200
rect 796 -1200 856 1200
<< ndiff >>
rect -914 1188 -856 1200
rect -914 -1188 -902 1188
rect -868 -1188 -856 1188
rect -914 -1200 -856 -1188
rect -796 1188 -738 1200
rect -796 -1188 -784 1188
rect -750 -1188 -738 1188
rect -796 -1200 -738 -1188
rect -678 1188 -620 1200
rect -678 -1188 -666 1188
rect -632 -1188 -620 1188
rect -678 -1200 -620 -1188
rect -560 1188 -502 1200
rect -560 -1188 -548 1188
rect -514 -1188 -502 1188
rect -560 -1200 -502 -1188
rect -442 1188 -384 1200
rect -442 -1188 -430 1188
rect -396 -1188 -384 1188
rect -442 -1200 -384 -1188
rect -324 1188 -266 1200
rect -324 -1188 -312 1188
rect -278 -1188 -266 1188
rect -324 -1200 -266 -1188
rect -206 1188 -148 1200
rect -206 -1188 -194 1188
rect -160 -1188 -148 1188
rect -206 -1200 -148 -1188
rect -88 1188 -30 1200
rect -88 -1188 -76 1188
rect -42 -1188 -30 1188
rect -88 -1200 -30 -1188
rect 30 1188 88 1200
rect 30 -1188 42 1188
rect 76 -1188 88 1188
rect 30 -1200 88 -1188
rect 148 1188 206 1200
rect 148 -1188 160 1188
rect 194 -1188 206 1188
rect 148 -1200 206 -1188
rect 266 1188 324 1200
rect 266 -1188 278 1188
rect 312 -1188 324 1188
rect 266 -1200 324 -1188
rect 384 1188 442 1200
rect 384 -1188 396 1188
rect 430 -1188 442 1188
rect 384 -1200 442 -1188
rect 502 1188 560 1200
rect 502 -1188 514 1188
rect 548 -1188 560 1188
rect 502 -1200 560 -1188
rect 620 1188 678 1200
rect 620 -1188 632 1188
rect 666 -1188 678 1188
rect 620 -1200 678 -1188
rect 738 1188 796 1200
rect 738 -1188 750 1188
rect 784 -1188 796 1188
rect 738 -1200 796 -1188
rect 856 1188 914 1200
rect 856 -1188 868 1188
rect 902 -1188 914 1188
rect 856 -1200 914 -1188
<< ndiffc >>
rect -902 -1188 -868 1188
rect -784 -1188 -750 1188
rect -666 -1188 -632 1188
rect -548 -1188 -514 1188
rect -430 -1188 -396 1188
rect -312 -1188 -278 1188
rect -194 -1188 -160 1188
rect -76 -1188 -42 1188
rect 42 -1188 76 1188
rect 160 -1188 194 1188
rect 278 -1188 312 1188
rect 396 -1188 430 1188
rect 514 -1188 548 1188
rect 632 -1188 666 1188
rect 750 -1188 784 1188
rect 868 -1188 902 1188
<< psubdiff >>
rect -1016 1340 -920 1374
rect 920 1340 1016 1374
rect -1016 1278 -982 1340
rect 982 1278 1016 1340
rect -1016 -1340 -982 -1278
rect 982 -1340 1016 -1278
rect -1016 -1374 -920 -1340
rect 920 -1374 1016 -1340
<< psubdiffcont >>
rect -920 1340 920 1374
rect -1016 -1278 -982 1278
rect 982 -1278 1016 1278
rect -920 -1374 920 -1340
<< poly >>
rect -859 1272 -793 1288
rect -859 1238 -843 1272
rect -809 1238 -793 1272
rect -859 1222 -793 1238
rect -741 1272 -675 1288
rect -741 1238 -725 1272
rect -691 1238 -675 1272
rect -741 1222 -675 1238
rect -623 1272 -557 1288
rect -623 1238 -607 1272
rect -573 1238 -557 1272
rect -623 1222 -557 1238
rect -505 1272 -439 1288
rect -505 1238 -489 1272
rect -455 1238 -439 1272
rect -505 1222 -439 1238
rect -387 1272 -321 1288
rect -387 1238 -371 1272
rect -337 1238 -321 1272
rect -387 1222 -321 1238
rect -269 1272 -203 1288
rect -269 1238 -253 1272
rect -219 1238 -203 1272
rect -269 1222 -203 1238
rect -151 1272 -85 1288
rect -151 1238 -135 1272
rect -101 1238 -85 1272
rect -151 1222 -85 1238
rect -33 1272 33 1288
rect -33 1238 -17 1272
rect 17 1238 33 1272
rect -33 1222 33 1238
rect 85 1272 151 1288
rect 85 1238 101 1272
rect 135 1238 151 1272
rect 85 1222 151 1238
rect 203 1272 269 1288
rect 203 1238 219 1272
rect 253 1238 269 1272
rect 203 1222 269 1238
rect 321 1272 387 1288
rect 321 1238 337 1272
rect 371 1238 387 1272
rect 321 1222 387 1238
rect 439 1272 505 1288
rect 439 1238 455 1272
rect 489 1238 505 1272
rect 439 1222 505 1238
rect 557 1272 623 1288
rect 557 1238 573 1272
rect 607 1238 623 1272
rect 557 1222 623 1238
rect 675 1272 741 1288
rect 675 1238 691 1272
rect 725 1238 741 1272
rect 675 1222 741 1238
rect 793 1272 859 1288
rect 793 1238 809 1272
rect 843 1238 859 1272
rect 793 1222 859 1238
rect -856 1200 -796 1222
rect -738 1200 -678 1222
rect -620 1200 -560 1222
rect -502 1200 -442 1222
rect -384 1200 -324 1222
rect -266 1200 -206 1222
rect -148 1200 -88 1222
rect -30 1200 30 1222
rect 88 1200 148 1222
rect 206 1200 266 1222
rect 324 1200 384 1222
rect 442 1200 502 1222
rect 560 1200 620 1222
rect 678 1200 738 1222
rect 796 1200 856 1222
rect -856 -1222 -796 -1200
rect -738 -1222 -678 -1200
rect -620 -1222 -560 -1200
rect -502 -1222 -442 -1200
rect -384 -1222 -324 -1200
rect -266 -1222 -206 -1200
rect -148 -1222 -88 -1200
rect -30 -1222 30 -1200
rect 88 -1222 148 -1200
rect 206 -1222 266 -1200
rect 324 -1222 384 -1200
rect 442 -1222 502 -1200
rect 560 -1222 620 -1200
rect 678 -1222 738 -1200
rect 796 -1222 856 -1200
rect -859 -1238 -793 -1222
rect -859 -1272 -843 -1238
rect -809 -1272 -793 -1238
rect -859 -1288 -793 -1272
rect -741 -1238 -675 -1222
rect -741 -1272 -725 -1238
rect -691 -1272 -675 -1238
rect -741 -1288 -675 -1272
rect -623 -1238 -557 -1222
rect -623 -1272 -607 -1238
rect -573 -1272 -557 -1238
rect -623 -1288 -557 -1272
rect -505 -1238 -439 -1222
rect -505 -1272 -489 -1238
rect -455 -1272 -439 -1238
rect -505 -1288 -439 -1272
rect -387 -1238 -321 -1222
rect -387 -1272 -371 -1238
rect -337 -1272 -321 -1238
rect -387 -1288 -321 -1272
rect -269 -1238 -203 -1222
rect -269 -1272 -253 -1238
rect -219 -1272 -203 -1238
rect -269 -1288 -203 -1272
rect -151 -1238 -85 -1222
rect -151 -1272 -135 -1238
rect -101 -1272 -85 -1238
rect -151 -1288 -85 -1272
rect -33 -1238 33 -1222
rect -33 -1272 -17 -1238
rect 17 -1272 33 -1238
rect -33 -1288 33 -1272
rect 85 -1238 151 -1222
rect 85 -1272 101 -1238
rect 135 -1272 151 -1238
rect 85 -1288 151 -1272
rect 203 -1238 269 -1222
rect 203 -1272 219 -1238
rect 253 -1272 269 -1238
rect 203 -1288 269 -1272
rect 321 -1238 387 -1222
rect 321 -1272 337 -1238
rect 371 -1272 387 -1238
rect 321 -1288 387 -1272
rect 439 -1238 505 -1222
rect 439 -1272 455 -1238
rect 489 -1272 505 -1238
rect 439 -1288 505 -1272
rect 557 -1238 623 -1222
rect 557 -1272 573 -1238
rect 607 -1272 623 -1238
rect 557 -1288 623 -1272
rect 675 -1238 741 -1222
rect 675 -1272 691 -1238
rect 725 -1272 741 -1238
rect 675 -1288 741 -1272
rect 793 -1238 859 -1222
rect 793 -1272 809 -1238
rect 843 -1272 859 -1238
rect 793 -1288 859 -1272
<< polycont >>
rect -843 1238 -809 1272
rect -725 1238 -691 1272
rect -607 1238 -573 1272
rect -489 1238 -455 1272
rect -371 1238 -337 1272
rect -253 1238 -219 1272
rect -135 1238 -101 1272
rect -17 1238 17 1272
rect 101 1238 135 1272
rect 219 1238 253 1272
rect 337 1238 371 1272
rect 455 1238 489 1272
rect 573 1238 607 1272
rect 691 1238 725 1272
rect 809 1238 843 1272
rect -843 -1272 -809 -1238
rect -725 -1272 -691 -1238
rect -607 -1272 -573 -1238
rect -489 -1272 -455 -1238
rect -371 -1272 -337 -1238
rect -253 -1272 -219 -1238
rect -135 -1272 -101 -1238
rect -17 -1272 17 -1238
rect 101 -1272 135 -1238
rect 219 -1272 253 -1238
rect 337 -1272 371 -1238
rect 455 -1272 489 -1238
rect 573 -1272 607 -1238
rect 691 -1272 725 -1238
rect 809 -1272 843 -1238
<< locali >>
rect -1016 1340 -920 1374
rect 920 1340 1016 1374
rect -1016 1278 -982 1340
rect 982 1278 1016 1340
rect -859 1238 -843 1272
rect -809 1238 -793 1272
rect -741 1238 -725 1272
rect -691 1238 -675 1272
rect -623 1238 -607 1272
rect -573 1238 -557 1272
rect -505 1238 -489 1272
rect -455 1238 -439 1272
rect -387 1238 -371 1272
rect -337 1238 -321 1272
rect -269 1238 -253 1272
rect -219 1238 -203 1272
rect -151 1238 -135 1272
rect -101 1238 -85 1272
rect -33 1238 -17 1272
rect 17 1238 33 1272
rect 85 1238 101 1272
rect 135 1238 151 1272
rect 203 1238 219 1272
rect 253 1238 269 1272
rect 321 1238 337 1272
rect 371 1238 387 1272
rect 439 1238 455 1272
rect 489 1238 505 1272
rect 557 1238 573 1272
rect 607 1238 623 1272
rect 675 1238 691 1272
rect 725 1238 741 1272
rect 793 1238 809 1272
rect 843 1238 859 1272
rect -902 1188 -868 1204
rect -902 -1204 -868 -1188
rect -784 1188 -750 1204
rect -784 -1204 -750 -1188
rect -666 1188 -632 1204
rect -666 -1204 -632 -1188
rect -548 1188 -514 1204
rect -548 -1204 -514 -1188
rect -430 1188 -396 1204
rect -430 -1204 -396 -1188
rect -312 1188 -278 1204
rect -312 -1204 -278 -1188
rect -194 1188 -160 1204
rect -194 -1204 -160 -1188
rect -76 1188 -42 1204
rect -76 -1204 -42 -1188
rect 42 1188 76 1204
rect 42 -1204 76 -1188
rect 160 1188 194 1204
rect 160 -1204 194 -1188
rect 278 1188 312 1204
rect 278 -1204 312 -1188
rect 396 1188 430 1204
rect 396 -1204 430 -1188
rect 514 1188 548 1204
rect 514 -1204 548 -1188
rect 632 1188 666 1204
rect 632 -1204 666 -1188
rect 750 1188 784 1204
rect 750 -1204 784 -1188
rect 868 1188 902 1204
rect 868 -1204 902 -1188
rect -859 -1272 -843 -1238
rect -809 -1272 -793 -1238
rect -741 -1272 -725 -1238
rect -691 -1272 -675 -1238
rect -623 -1272 -607 -1238
rect -573 -1272 -557 -1238
rect -505 -1272 -489 -1238
rect -455 -1272 -439 -1238
rect -387 -1272 -371 -1238
rect -337 -1272 -321 -1238
rect -269 -1272 -253 -1238
rect -219 -1272 -203 -1238
rect -151 -1272 -135 -1238
rect -101 -1272 -85 -1238
rect -33 -1272 -17 -1238
rect 17 -1272 33 -1238
rect 85 -1272 101 -1238
rect 135 -1272 151 -1238
rect 203 -1272 219 -1238
rect 253 -1272 269 -1238
rect 321 -1272 337 -1238
rect 371 -1272 387 -1238
rect 439 -1272 455 -1238
rect 489 -1272 505 -1238
rect 557 -1272 573 -1238
rect 607 -1272 623 -1238
rect 675 -1272 691 -1238
rect 725 -1272 741 -1238
rect 793 -1272 809 -1238
rect 843 -1272 859 -1238
rect -1016 -1340 -982 -1278
rect 982 -1340 1016 -1278
rect -1016 -1374 -920 -1340
rect 920 -1374 1016 -1340
<< viali >>
rect -843 1238 -809 1272
rect -725 1238 -691 1272
rect -607 1238 -573 1272
rect -489 1238 -455 1272
rect -371 1238 -337 1272
rect -253 1238 -219 1272
rect -135 1238 -101 1272
rect -17 1238 17 1272
rect 101 1238 135 1272
rect 219 1238 253 1272
rect 337 1238 371 1272
rect 455 1238 489 1272
rect 573 1238 607 1272
rect 691 1238 725 1272
rect 809 1238 843 1272
rect -902 -1188 -868 1188
rect -784 -1188 -750 1188
rect -666 -1188 -632 1188
rect -548 -1188 -514 1188
rect -430 -1188 -396 1188
rect -312 -1188 -278 1188
rect -194 -1188 -160 1188
rect -76 -1188 -42 1188
rect 42 -1188 76 1188
rect 160 -1188 194 1188
rect 278 -1188 312 1188
rect 396 -1188 430 1188
rect 514 -1188 548 1188
rect 632 -1188 666 1188
rect 750 -1188 784 1188
rect 868 -1188 902 1188
rect -843 -1272 -809 -1238
rect -725 -1272 -691 -1238
rect -607 -1272 -573 -1238
rect -489 -1272 -455 -1238
rect -371 -1272 -337 -1238
rect -253 -1272 -219 -1238
rect -135 -1272 -101 -1238
rect -17 -1272 17 -1238
rect 101 -1272 135 -1238
rect 219 -1272 253 -1238
rect 337 -1272 371 -1238
rect 455 -1272 489 -1238
rect 573 -1272 607 -1238
rect 691 -1272 725 -1238
rect 809 -1272 843 -1238
<< metal1 >>
rect -855 1272 -797 1278
rect -855 1238 -843 1272
rect -809 1238 -797 1272
rect -855 1232 -797 1238
rect -737 1272 -679 1278
rect -737 1238 -725 1272
rect -691 1238 -679 1272
rect -737 1232 -679 1238
rect -619 1272 -561 1278
rect -619 1238 -607 1272
rect -573 1238 -561 1272
rect -619 1232 -561 1238
rect -501 1272 -443 1278
rect -501 1238 -489 1272
rect -455 1238 -443 1272
rect -501 1232 -443 1238
rect -383 1272 -325 1278
rect -383 1238 -371 1272
rect -337 1238 -325 1272
rect -383 1232 -325 1238
rect -265 1272 -207 1278
rect -265 1238 -253 1272
rect -219 1238 -207 1272
rect -265 1232 -207 1238
rect -147 1272 -89 1278
rect -147 1238 -135 1272
rect -101 1238 -89 1272
rect -147 1232 -89 1238
rect -29 1272 29 1278
rect -29 1238 -17 1272
rect 17 1238 29 1272
rect -29 1232 29 1238
rect 89 1272 147 1278
rect 89 1238 101 1272
rect 135 1238 147 1272
rect 89 1232 147 1238
rect 207 1272 265 1278
rect 207 1238 219 1272
rect 253 1238 265 1272
rect 207 1232 265 1238
rect 325 1272 383 1278
rect 325 1238 337 1272
rect 371 1238 383 1272
rect 325 1232 383 1238
rect 443 1272 501 1278
rect 443 1238 455 1272
rect 489 1238 501 1272
rect 443 1232 501 1238
rect 561 1272 619 1278
rect 561 1238 573 1272
rect 607 1238 619 1272
rect 561 1232 619 1238
rect 679 1272 737 1278
rect 679 1238 691 1272
rect 725 1238 737 1272
rect 679 1232 737 1238
rect 797 1272 855 1278
rect 797 1238 809 1272
rect 843 1238 855 1272
rect 797 1232 855 1238
rect -908 1188 -862 1200
rect -908 -1188 -902 1188
rect -868 -1188 -862 1188
rect -908 -1200 -862 -1188
rect -790 1188 -744 1200
rect -790 -1188 -784 1188
rect -750 -1188 -744 1188
rect -790 -1200 -744 -1188
rect -672 1188 -626 1200
rect -672 -1188 -666 1188
rect -632 -1188 -626 1188
rect -672 -1200 -626 -1188
rect -554 1188 -508 1200
rect -554 -1188 -548 1188
rect -514 -1188 -508 1188
rect -554 -1200 -508 -1188
rect -436 1188 -390 1200
rect -436 -1188 -430 1188
rect -396 -1188 -390 1188
rect -436 -1200 -390 -1188
rect -318 1188 -272 1200
rect -318 -1188 -312 1188
rect -278 -1188 -272 1188
rect -318 -1200 -272 -1188
rect -200 1188 -154 1200
rect -200 -1188 -194 1188
rect -160 -1188 -154 1188
rect -200 -1200 -154 -1188
rect -82 1188 -36 1200
rect -82 -1188 -76 1188
rect -42 -1188 -36 1188
rect -82 -1200 -36 -1188
rect 36 1188 82 1200
rect 36 -1188 42 1188
rect 76 -1188 82 1188
rect 36 -1200 82 -1188
rect 154 1188 200 1200
rect 154 -1188 160 1188
rect 194 -1188 200 1188
rect 154 -1200 200 -1188
rect 272 1188 318 1200
rect 272 -1188 278 1188
rect 312 -1188 318 1188
rect 272 -1200 318 -1188
rect 390 1188 436 1200
rect 390 -1188 396 1188
rect 430 -1188 436 1188
rect 390 -1200 436 -1188
rect 508 1188 554 1200
rect 508 -1188 514 1188
rect 548 -1188 554 1188
rect 508 -1200 554 -1188
rect 626 1188 672 1200
rect 626 -1188 632 1188
rect 666 -1188 672 1188
rect 626 -1200 672 -1188
rect 744 1188 790 1200
rect 744 -1188 750 1188
rect 784 -1188 790 1188
rect 744 -1200 790 -1188
rect 862 1188 908 1200
rect 862 -1188 868 1188
rect 902 -1188 908 1188
rect 862 -1200 908 -1188
rect -855 -1238 -797 -1232
rect -855 -1272 -843 -1238
rect -809 -1272 -797 -1238
rect -855 -1278 -797 -1272
rect -737 -1238 -679 -1232
rect -737 -1272 -725 -1238
rect -691 -1272 -679 -1238
rect -737 -1278 -679 -1272
rect -619 -1238 -561 -1232
rect -619 -1272 -607 -1238
rect -573 -1272 -561 -1238
rect -619 -1278 -561 -1272
rect -501 -1238 -443 -1232
rect -501 -1272 -489 -1238
rect -455 -1272 -443 -1238
rect -501 -1278 -443 -1272
rect -383 -1238 -325 -1232
rect -383 -1272 -371 -1238
rect -337 -1272 -325 -1238
rect -383 -1278 -325 -1272
rect -265 -1238 -207 -1232
rect -265 -1272 -253 -1238
rect -219 -1272 -207 -1238
rect -265 -1278 -207 -1272
rect -147 -1238 -89 -1232
rect -147 -1272 -135 -1238
rect -101 -1272 -89 -1238
rect -147 -1278 -89 -1272
rect -29 -1238 29 -1232
rect -29 -1272 -17 -1238
rect 17 -1272 29 -1238
rect -29 -1278 29 -1272
rect 89 -1238 147 -1232
rect 89 -1272 101 -1238
rect 135 -1272 147 -1238
rect 89 -1278 147 -1272
rect 207 -1238 265 -1232
rect 207 -1272 219 -1238
rect 253 -1272 265 -1238
rect 207 -1278 265 -1272
rect 325 -1238 383 -1232
rect 325 -1272 337 -1238
rect 371 -1272 383 -1238
rect 325 -1278 383 -1272
rect 443 -1238 501 -1232
rect 443 -1272 455 -1238
rect 489 -1272 501 -1238
rect 443 -1278 501 -1272
rect 561 -1238 619 -1232
rect 561 -1272 573 -1238
rect 607 -1272 619 -1238
rect 561 -1278 619 -1272
rect 679 -1238 737 -1232
rect 679 -1272 691 -1238
rect 725 -1272 737 -1238
rect 679 -1278 737 -1272
rect 797 -1238 855 -1232
rect 797 -1272 809 -1238
rect 843 -1272 855 -1238
rect 797 -1278 855 -1272
<< properties >>
string FIXED_BBOX -999 -1357 999 1357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 12 l 0.30 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
