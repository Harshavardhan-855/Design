magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -125 1881 -67 1887
rect 67 1881 125 1887
rect -125 1847 -113 1881
rect 67 1847 79 1881
rect -125 1841 -67 1847
rect 67 1841 125 1847
rect -221 -1847 -163 -1841
rect -29 -1847 29 -1841
rect 163 -1847 221 -1841
rect -221 -1881 -209 -1847
rect -29 -1881 -17 -1847
rect 163 -1881 175 -1847
rect -221 -1887 -163 -1881
rect -29 -1887 29 -1881
rect 163 -1887 221 -1881
<< nwell >>
rect -407 -2019 407 2019
<< pmos >>
rect -207 -1800 -177 1800
rect -111 -1800 -81 1800
rect -15 -1800 15 1800
rect 81 -1800 111 1800
rect 177 -1800 207 1800
<< pdiff >>
rect -269 1788 -207 1800
rect -269 -1788 -257 1788
rect -223 -1788 -207 1788
rect -269 -1800 -207 -1788
rect -177 1788 -111 1800
rect -177 -1788 -161 1788
rect -127 -1788 -111 1788
rect -177 -1800 -111 -1788
rect -81 1788 -15 1800
rect -81 -1788 -65 1788
rect -31 -1788 -15 1788
rect -81 -1800 -15 -1788
rect 15 1788 81 1800
rect 15 -1788 31 1788
rect 65 -1788 81 1788
rect 15 -1800 81 -1788
rect 111 1788 177 1800
rect 111 -1788 127 1788
rect 161 -1788 177 1788
rect 111 -1800 177 -1788
rect 207 1788 269 1800
rect 207 -1788 223 1788
rect 257 -1788 269 1788
rect 207 -1800 269 -1788
<< pdiffc >>
rect -257 -1788 -223 1788
rect -161 -1788 -127 1788
rect -65 -1788 -31 1788
rect 31 -1788 65 1788
rect 127 -1788 161 1788
rect 223 -1788 257 1788
<< nsubdiff >>
rect -371 1949 -275 1983
rect 275 1949 371 1983
rect -371 1887 -337 1949
rect 337 1887 371 1949
rect -371 -1949 -337 -1887
rect 337 -1949 371 -1887
rect -371 -1983 -275 -1949
rect 275 -1983 371 -1949
<< nsubdiffcont >>
rect -275 1949 275 1983
rect -371 -1887 -337 1887
rect 337 -1887 371 1887
rect -275 -1983 275 -1949
<< poly >>
rect -129 1881 -63 1897
rect -129 1847 -113 1881
rect -79 1847 -63 1881
rect -129 1831 -63 1847
rect 63 1881 129 1897
rect 63 1847 79 1881
rect 113 1847 129 1881
rect 63 1831 129 1847
rect -207 1800 -177 1826
rect -111 1800 -81 1831
rect -15 1800 15 1826
rect 81 1800 111 1831
rect 177 1800 207 1826
rect -207 -1831 -177 -1800
rect -111 -1826 -81 -1800
rect -15 -1831 15 -1800
rect 81 -1826 111 -1800
rect 177 -1831 207 -1800
rect -225 -1847 -159 -1831
rect -225 -1881 -209 -1847
rect -175 -1881 -159 -1847
rect -225 -1897 -159 -1881
rect -33 -1847 33 -1831
rect -33 -1881 -17 -1847
rect 17 -1881 33 -1847
rect -33 -1897 33 -1881
rect 159 -1847 225 -1831
rect 159 -1881 175 -1847
rect 209 -1881 225 -1847
rect 159 -1897 225 -1881
<< polycont >>
rect -113 1847 -79 1881
rect 79 1847 113 1881
rect -209 -1881 -175 -1847
rect -17 -1881 17 -1847
rect 175 -1881 209 -1847
<< locali >>
rect -371 1949 -275 1983
rect 275 1949 371 1983
rect -371 1887 -337 1949
rect 337 1887 371 1949
rect -129 1847 -113 1881
rect -79 1847 -63 1881
rect 63 1847 79 1881
rect 113 1847 129 1881
rect -257 1788 -223 1804
rect -257 -1804 -223 -1788
rect -161 1788 -127 1804
rect -161 -1804 -127 -1788
rect -65 1788 -31 1804
rect -65 -1804 -31 -1788
rect 31 1788 65 1804
rect 31 -1804 65 -1788
rect 127 1788 161 1804
rect 127 -1804 161 -1788
rect 223 1788 257 1804
rect 223 -1804 257 -1788
rect -225 -1881 -209 -1847
rect -175 -1881 -159 -1847
rect -33 -1881 -17 -1847
rect 17 -1881 33 -1847
rect 159 -1881 175 -1847
rect 209 -1881 225 -1847
rect -371 -1949 -337 -1887
rect 337 -1949 371 -1887
rect -371 -1983 -275 -1949
rect 275 -1983 371 -1949
<< viali >>
rect -113 1847 -79 1881
rect 79 1847 113 1881
rect -257 -1788 -223 1788
rect -161 -1788 -127 1788
rect -65 -1788 -31 1788
rect 31 -1788 65 1788
rect 127 -1788 161 1788
rect 223 -1788 257 1788
rect -209 -1881 -175 -1847
rect -17 -1881 17 -1847
rect 175 -1881 209 -1847
<< metal1 >>
rect -125 1881 -67 1887
rect -125 1847 -113 1881
rect -79 1847 -67 1881
rect -125 1841 -67 1847
rect 67 1881 125 1887
rect 67 1847 79 1881
rect 113 1847 125 1881
rect 67 1841 125 1847
rect -263 1788 -217 1800
rect -263 -1788 -257 1788
rect -223 -1788 -217 1788
rect -263 -1800 -217 -1788
rect -167 1788 -121 1800
rect -167 -1788 -161 1788
rect -127 -1788 -121 1788
rect -167 -1800 -121 -1788
rect -71 1788 -25 1800
rect -71 -1788 -65 1788
rect -31 -1788 -25 1788
rect -71 -1800 -25 -1788
rect 25 1788 71 1800
rect 25 -1788 31 1788
rect 65 -1788 71 1788
rect 25 -1800 71 -1788
rect 121 1788 167 1800
rect 121 -1788 127 1788
rect 161 -1788 167 1788
rect 121 -1800 167 -1788
rect 217 1788 263 1800
rect 217 -1788 223 1788
rect 257 -1788 263 1788
rect 217 -1800 263 -1788
rect -221 -1847 -163 -1841
rect -221 -1881 -209 -1847
rect -175 -1881 -163 -1847
rect -221 -1887 -163 -1881
rect -29 -1847 29 -1841
rect -29 -1881 -17 -1847
rect 17 -1881 29 -1847
rect -29 -1887 29 -1881
rect 163 -1847 221 -1841
rect 163 -1881 175 -1847
rect 209 -1881 221 -1847
rect 163 -1887 221 -1881
<< properties >>
string FIXED_BBOX -354 -1966 354 1966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 18 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
