magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -845 881 -787 887
rect -653 881 -595 887
rect -461 881 -403 887
rect -269 881 -211 887
rect -77 881 -19 887
rect 115 881 173 887
rect 307 881 365 887
rect 499 881 557 887
rect 691 881 749 887
rect 883 881 941 887
rect -845 847 -833 881
rect -653 847 -641 881
rect -461 847 -449 881
rect -269 847 -257 881
rect -77 847 -65 881
rect 115 847 127 881
rect 307 847 319 881
rect 499 847 511 881
rect 691 847 703 881
rect 883 847 895 881
rect -845 841 -787 847
rect -653 841 -595 847
rect -461 841 -403 847
rect -269 841 -211 847
rect -77 841 -19 847
rect 115 841 173 847
rect 307 841 365 847
rect 499 841 557 847
rect 691 841 749 847
rect 883 841 941 847
rect -941 -847 -883 -841
rect -749 -847 -691 -841
rect -557 -847 -499 -841
rect -365 -847 -307 -841
rect -173 -847 -115 -841
rect 19 -847 77 -841
rect 211 -847 269 -841
rect 403 -847 461 -841
rect 595 -847 653 -841
rect 787 -847 845 -841
rect -941 -881 -929 -847
rect -749 -881 -737 -847
rect -557 -881 -545 -847
rect -365 -881 -353 -847
rect -173 -881 -161 -847
rect 19 -881 31 -847
rect 211 -881 223 -847
rect 403 -881 415 -847
rect 595 -881 607 -847
rect 787 -881 799 -847
rect -941 -887 -883 -881
rect -749 -887 -691 -881
rect -557 -887 -499 -881
rect -365 -887 -307 -881
rect -173 -887 -115 -881
rect 19 -887 77 -881
rect 211 -887 269 -881
rect 403 -887 461 -881
rect 595 -887 653 -881
rect 787 -887 845 -881
<< nwell >>
rect -1127 -1019 1127 1019
<< pmos >>
rect -927 -800 -897 800
rect -831 -800 -801 800
rect -735 -800 -705 800
rect -639 -800 -609 800
rect -543 -800 -513 800
rect -447 -800 -417 800
rect -351 -800 -321 800
rect -255 -800 -225 800
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
rect 225 -800 255 800
rect 321 -800 351 800
rect 417 -800 447 800
rect 513 -800 543 800
rect 609 -800 639 800
rect 705 -800 735 800
rect 801 -800 831 800
rect 897 -800 927 800
<< pdiff >>
rect -989 788 -927 800
rect -989 -788 -977 788
rect -943 -788 -927 788
rect -989 -800 -927 -788
rect -897 788 -831 800
rect -897 -788 -881 788
rect -847 -788 -831 788
rect -897 -800 -831 -788
rect -801 788 -735 800
rect -801 -788 -785 788
rect -751 -788 -735 788
rect -801 -800 -735 -788
rect -705 788 -639 800
rect -705 -788 -689 788
rect -655 -788 -639 788
rect -705 -800 -639 -788
rect -609 788 -543 800
rect -609 -788 -593 788
rect -559 -788 -543 788
rect -609 -800 -543 -788
rect -513 788 -447 800
rect -513 -788 -497 788
rect -463 -788 -447 788
rect -513 -800 -447 -788
rect -417 788 -351 800
rect -417 -788 -401 788
rect -367 -788 -351 788
rect -417 -800 -351 -788
rect -321 788 -255 800
rect -321 -788 -305 788
rect -271 -788 -255 788
rect -321 -800 -255 -788
rect -225 788 -159 800
rect -225 -788 -209 788
rect -175 -788 -159 788
rect -225 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 225 800
rect 159 -788 175 788
rect 209 -788 225 788
rect 159 -800 225 -788
rect 255 788 321 800
rect 255 -788 271 788
rect 305 -788 321 788
rect 255 -800 321 -788
rect 351 788 417 800
rect 351 -788 367 788
rect 401 -788 417 788
rect 351 -800 417 -788
rect 447 788 513 800
rect 447 -788 463 788
rect 497 -788 513 788
rect 447 -800 513 -788
rect 543 788 609 800
rect 543 -788 559 788
rect 593 -788 609 788
rect 543 -800 609 -788
rect 639 788 705 800
rect 639 -788 655 788
rect 689 -788 705 788
rect 639 -800 705 -788
rect 735 788 801 800
rect 735 -788 751 788
rect 785 -788 801 788
rect 735 -800 801 -788
rect 831 788 897 800
rect 831 -788 847 788
rect 881 -788 897 788
rect 831 -800 897 -788
rect 927 788 989 800
rect 927 -788 943 788
rect 977 -788 989 788
rect 927 -800 989 -788
<< pdiffc >>
rect -977 -788 -943 788
rect -881 -788 -847 788
rect -785 -788 -751 788
rect -689 -788 -655 788
rect -593 -788 -559 788
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect 559 -788 593 788
rect 655 -788 689 788
rect 751 -788 785 788
rect 847 -788 881 788
rect 943 -788 977 788
<< nsubdiff >>
rect -1091 949 -995 983
rect 995 949 1091 983
rect -1091 887 -1057 949
rect 1057 887 1091 949
rect -1091 -949 -1057 -887
rect 1057 -949 1091 -887
rect -1091 -983 -995 -949
rect 995 -983 1091 -949
<< nsubdiffcont >>
rect -995 949 995 983
rect -1091 -887 -1057 887
rect 1057 -887 1091 887
rect -995 -983 995 -949
<< poly >>
rect -849 881 -783 897
rect -849 847 -833 881
rect -799 847 -783 881
rect -849 831 -783 847
rect -657 881 -591 897
rect -657 847 -641 881
rect -607 847 -591 881
rect -657 831 -591 847
rect -465 881 -399 897
rect -465 847 -449 881
rect -415 847 -399 881
rect -465 831 -399 847
rect -273 881 -207 897
rect -273 847 -257 881
rect -223 847 -207 881
rect -273 831 -207 847
rect -81 881 -15 897
rect -81 847 -65 881
rect -31 847 -15 881
rect -81 831 -15 847
rect 111 881 177 897
rect 111 847 127 881
rect 161 847 177 881
rect 111 831 177 847
rect 303 881 369 897
rect 303 847 319 881
rect 353 847 369 881
rect 303 831 369 847
rect 495 881 561 897
rect 495 847 511 881
rect 545 847 561 881
rect 495 831 561 847
rect 687 881 753 897
rect 687 847 703 881
rect 737 847 753 881
rect 687 831 753 847
rect 879 881 945 897
rect 879 847 895 881
rect 929 847 945 881
rect 879 831 945 847
rect -927 800 -897 826
rect -831 800 -801 831
rect -735 800 -705 826
rect -639 800 -609 831
rect -543 800 -513 826
rect -447 800 -417 831
rect -351 800 -321 826
rect -255 800 -225 831
rect -159 800 -129 826
rect -63 800 -33 831
rect 33 800 63 826
rect 129 800 159 831
rect 225 800 255 826
rect 321 800 351 831
rect 417 800 447 826
rect 513 800 543 831
rect 609 800 639 826
rect 705 800 735 831
rect 801 800 831 826
rect 897 800 927 831
rect -927 -831 -897 -800
rect -831 -826 -801 -800
rect -735 -831 -705 -800
rect -639 -826 -609 -800
rect -543 -831 -513 -800
rect -447 -826 -417 -800
rect -351 -831 -321 -800
rect -255 -826 -225 -800
rect -159 -831 -129 -800
rect -63 -826 -33 -800
rect 33 -831 63 -800
rect 129 -826 159 -800
rect 225 -831 255 -800
rect 321 -826 351 -800
rect 417 -831 447 -800
rect 513 -826 543 -800
rect 609 -831 639 -800
rect 705 -826 735 -800
rect 801 -831 831 -800
rect 897 -826 927 -800
rect -945 -847 -879 -831
rect -945 -881 -929 -847
rect -895 -881 -879 -847
rect -945 -897 -879 -881
rect -753 -847 -687 -831
rect -753 -881 -737 -847
rect -703 -881 -687 -847
rect -753 -897 -687 -881
rect -561 -847 -495 -831
rect -561 -881 -545 -847
rect -511 -881 -495 -847
rect -561 -897 -495 -881
rect -369 -847 -303 -831
rect -369 -881 -353 -847
rect -319 -881 -303 -847
rect -369 -897 -303 -881
rect -177 -847 -111 -831
rect -177 -881 -161 -847
rect -127 -881 -111 -847
rect -177 -897 -111 -881
rect 15 -847 81 -831
rect 15 -881 31 -847
rect 65 -881 81 -847
rect 15 -897 81 -881
rect 207 -847 273 -831
rect 207 -881 223 -847
rect 257 -881 273 -847
rect 207 -897 273 -881
rect 399 -847 465 -831
rect 399 -881 415 -847
rect 449 -881 465 -847
rect 399 -897 465 -881
rect 591 -847 657 -831
rect 591 -881 607 -847
rect 641 -881 657 -847
rect 591 -897 657 -881
rect 783 -847 849 -831
rect 783 -881 799 -847
rect 833 -881 849 -847
rect 783 -897 849 -881
<< polycont >>
rect -833 847 -799 881
rect -641 847 -607 881
rect -449 847 -415 881
rect -257 847 -223 881
rect -65 847 -31 881
rect 127 847 161 881
rect 319 847 353 881
rect 511 847 545 881
rect 703 847 737 881
rect 895 847 929 881
rect -929 -881 -895 -847
rect -737 -881 -703 -847
rect -545 -881 -511 -847
rect -353 -881 -319 -847
rect -161 -881 -127 -847
rect 31 -881 65 -847
rect 223 -881 257 -847
rect 415 -881 449 -847
rect 607 -881 641 -847
rect 799 -881 833 -847
<< locali >>
rect -1091 949 -995 983
rect 995 949 1091 983
rect -1091 887 -1057 949
rect 1057 887 1091 949
rect -849 847 -833 881
rect -799 847 -783 881
rect -657 847 -641 881
rect -607 847 -591 881
rect -465 847 -449 881
rect -415 847 -399 881
rect -273 847 -257 881
rect -223 847 -207 881
rect -81 847 -65 881
rect -31 847 -15 881
rect 111 847 127 881
rect 161 847 177 881
rect 303 847 319 881
rect 353 847 369 881
rect 495 847 511 881
rect 545 847 561 881
rect 687 847 703 881
rect 737 847 753 881
rect 879 847 895 881
rect 929 847 945 881
rect -977 788 -943 804
rect -977 -804 -943 -788
rect -881 788 -847 804
rect -881 -804 -847 -788
rect -785 788 -751 804
rect -785 -804 -751 -788
rect -689 788 -655 804
rect -689 -804 -655 -788
rect -593 788 -559 804
rect -593 -804 -559 -788
rect -497 788 -463 804
rect -497 -804 -463 -788
rect -401 788 -367 804
rect -401 -804 -367 -788
rect -305 788 -271 804
rect -305 -804 -271 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 271 788 305 804
rect 271 -804 305 -788
rect 367 788 401 804
rect 367 -804 401 -788
rect 463 788 497 804
rect 463 -804 497 -788
rect 559 788 593 804
rect 559 -804 593 -788
rect 655 788 689 804
rect 655 -804 689 -788
rect 751 788 785 804
rect 751 -804 785 -788
rect 847 788 881 804
rect 847 -804 881 -788
rect 943 788 977 804
rect 943 -804 977 -788
rect -945 -881 -929 -847
rect -895 -881 -879 -847
rect -753 -881 -737 -847
rect -703 -881 -687 -847
rect -561 -881 -545 -847
rect -511 -881 -495 -847
rect -369 -881 -353 -847
rect -319 -881 -303 -847
rect -177 -881 -161 -847
rect -127 -881 -111 -847
rect 15 -881 31 -847
rect 65 -881 81 -847
rect 207 -881 223 -847
rect 257 -881 273 -847
rect 399 -881 415 -847
rect 449 -881 465 -847
rect 591 -881 607 -847
rect 641 -881 657 -847
rect 783 -881 799 -847
rect 833 -881 849 -847
rect -1091 -949 -1057 -887
rect 1057 -949 1091 -887
rect -1091 -983 -995 -949
rect 995 -983 1091 -949
<< viali >>
rect -833 847 -799 881
rect -641 847 -607 881
rect -449 847 -415 881
rect -257 847 -223 881
rect -65 847 -31 881
rect 127 847 161 881
rect 319 847 353 881
rect 511 847 545 881
rect 703 847 737 881
rect 895 847 929 881
rect -977 -788 -943 788
rect -881 -788 -847 788
rect -785 -788 -751 788
rect -689 -788 -655 788
rect -593 -788 -559 788
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect 559 -788 593 788
rect 655 -788 689 788
rect 751 -788 785 788
rect 847 -788 881 788
rect 943 -788 977 788
rect -929 -881 -895 -847
rect -737 -881 -703 -847
rect -545 -881 -511 -847
rect -353 -881 -319 -847
rect -161 -881 -127 -847
rect 31 -881 65 -847
rect 223 -881 257 -847
rect 415 -881 449 -847
rect 607 -881 641 -847
rect 799 -881 833 -847
<< metal1 >>
rect -845 881 -787 887
rect -845 847 -833 881
rect -799 847 -787 881
rect -845 841 -787 847
rect -653 881 -595 887
rect -653 847 -641 881
rect -607 847 -595 881
rect -653 841 -595 847
rect -461 881 -403 887
rect -461 847 -449 881
rect -415 847 -403 881
rect -461 841 -403 847
rect -269 881 -211 887
rect -269 847 -257 881
rect -223 847 -211 881
rect -269 841 -211 847
rect -77 881 -19 887
rect -77 847 -65 881
rect -31 847 -19 881
rect -77 841 -19 847
rect 115 881 173 887
rect 115 847 127 881
rect 161 847 173 881
rect 115 841 173 847
rect 307 881 365 887
rect 307 847 319 881
rect 353 847 365 881
rect 307 841 365 847
rect 499 881 557 887
rect 499 847 511 881
rect 545 847 557 881
rect 499 841 557 847
rect 691 881 749 887
rect 691 847 703 881
rect 737 847 749 881
rect 691 841 749 847
rect 883 881 941 887
rect 883 847 895 881
rect 929 847 941 881
rect 883 841 941 847
rect -983 788 -937 800
rect -983 -788 -977 788
rect -943 -788 -937 788
rect -983 -800 -937 -788
rect -887 788 -841 800
rect -887 -788 -881 788
rect -847 -788 -841 788
rect -887 -800 -841 -788
rect -791 788 -745 800
rect -791 -788 -785 788
rect -751 -788 -745 788
rect -791 -800 -745 -788
rect -695 788 -649 800
rect -695 -788 -689 788
rect -655 -788 -649 788
rect -695 -800 -649 -788
rect -599 788 -553 800
rect -599 -788 -593 788
rect -559 -788 -553 788
rect -599 -800 -553 -788
rect -503 788 -457 800
rect -503 -788 -497 788
rect -463 -788 -457 788
rect -503 -800 -457 -788
rect -407 788 -361 800
rect -407 -788 -401 788
rect -367 -788 -361 788
rect -407 -800 -361 -788
rect -311 788 -265 800
rect -311 -788 -305 788
rect -271 -788 -265 788
rect -311 -800 -265 -788
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect 265 788 311 800
rect 265 -788 271 788
rect 305 -788 311 788
rect 265 -800 311 -788
rect 361 788 407 800
rect 361 -788 367 788
rect 401 -788 407 788
rect 361 -800 407 -788
rect 457 788 503 800
rect 457 -788 463 788
rect 497 -788 503 788
rect 457 -800 503 -788
rect 553 788 599 800
rect 553 -788 559 788
rect 593 -788 599 788
rect 553 -800 599 -788
rect 649 788 695 800
rect 649 -788 655 788
rect 689 -788 695 788
rect 649 -800 695 -788
rect 745 788 791 800
rect 745 -788 751 788
rect 785 -788 791 788
rect 745 -800 791 -788
rect 841 788 887 800
rect 841 -788 847 788
rect 881 -788 887 788
rect 841 -800 887 -788
rect 937 788 983 800
rect 937 -788 943 788
rect 977 -788 983 788
rect 937 -800 983 -788
rect -941 -847 -883 -841
rect -941 -881 -929 -847
rect -895 -881 -883 -847
rect -941 -887 -883 -881
rect -749 -847 -691 -841
rect -749 -881 -737 -847
rect -703 -881 -691 -847
rect -749 -887 -691 -881
rect -557 -847 -499 -841
rect -557 -881 -545 -847
rect -511 -881 -499 -847
rect -557 -887 -499 -881
rect -365 -847 -307 -841
rect -365 -881 -353 -847
rect -319 -881 -307 -847
rect -365 -887 -307 -881
rect -173 -847 -115 -841
rect -173 -881 -161 -847
rect -127 -881 -115 -847
rect -173 -887 -115 -881
rect 19 -847 77 -841
rect 19 -881 31 -847
rect 65 -881 77 -847
rect 19 -887 77 -881
rect 211 -847 269 -841
rect 211 -881 223 -847
rect 257 -881 269 -847
rect 211 -887 269 -881
rect 403 -847 461 -841
rect 403 -881 415 -847
rect 449 -881 461 -847
rect 403 -887 461 -881
rect 595 -847 653 -841
rect 595 -881 607 -847
rect 641 -881 653 -847
rect 595 -887 653 -881
rect 787 -847 845 -841
rect 787 -881 799 -847
rect 833 -881 845 -847
rect 787 -887 845 -881
<< properties >>
string FIXED_BBOX -1074 -966 1074 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
