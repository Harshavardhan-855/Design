magic
tech sky130A
timestamp 1709275732
<< end >>
