magic
tech sky130A
magscale 1 2
timestamp 1709276291
<< nwell >>
rect 3324 5556 3370 5558
rect 4758 5556 4804 5558
rect 1938 5522 4804 5556
rect 3324 5332 3370 5522
rect 4758 5332 4804 5522
rect 2192 5034 2450 5070
rect 2414 4826 2450 5034
rect 2414 4790 2692 4826
<< locali >>
rect 2604 5408 2672 5558
rect 4040 5406 4108 5556
rect 5468 5408 5536 5558
rect 2096 5068 2176 5216
rect 2776 4944 2884 5222
rect 5348 4950 5456 5228
rect 3774 4120 3904 4154
rect 4092 4116 4138 4264
rect 4674 4114 4720 4262
rect 5396 4118 5442 4266
<< viali >>
rect 1842 5422 1882 5460
rect 5746 4118 5788 4154
<< metal1 >>
rect 1302 5466 1502 5610
rect 3324 5552 3370 5554
rect 4758 5552 4804 5554
rect 6142 5552 6188 5554
rect 1938 5518 6188 5552
rect 1302 5460 1894 5466
rect 1302 5422 1842 5460
rect 1882 5422 1894 5460
rect 1302 5416 1894 5422
rect 1302 5410 1892 5416
rect 1938 5328 1992 5518
rect 3324 5398 3370 5518
rect 4758 5398 4804 5518
rect 3272 5330 3426 5398
rect 1488 5088 1626 5090
rect 1942 5088 1988 5328
rect 4702 5326 4864 5398
rect 6142 5328 6188 5518
rect 3208 5282 3236 5312
rect 3458 5282 3486 5312
rect 3208 5254 3486 5282
rect 4630 5292 4664 5304
rect 4902 5292 4936 5308
rect 4630 5262 4666 5292
rect 4900 5262 4936 5292
rect 4630 5234 4936 5262
rect 1298 5042 1988 5088
rect 1298 4888 1498 5042
rect 2192 5034 2450 5070
rect 2192 4950 2228 5034
rect 2414 4826 2450 5034
rect 2562 4882 2618 4950
rect 4094 4886 4346 4946
rect 2652 4826 2692 4874
rect 2414 4790 2692 4826
rect 4202 4762 4272 4886
rect 5624 4882 5680 4950
rect 4510 4762 4570 4878
rect 4202 4724 4570 4762
rect 4204 4706 4570 4724
rect 1302 4552 1990 4604
rect 2378 4588 2388 4682
rect 2474 4588 2484 4682
rect 1302 4404 1502 4552
rect 2162 4400 2206 4538
rect 2406 4400 2450 4588
rect 3674 4426 4132 4458
rect 2162 4356 2638 4400
rect 4094 4352 4132 4426
rect 4510 4350 4570 4706
rect 5836 4454 5904 5322
rect 6124 4706 6324 4748
rect 6124 4582 6178 4706
rect 6272 4582 6324 4706
rect 6124 4548 6324 4582
rect 5564 4422 5904 4454
rect 5564 4350 5612 4422
rect 3966 4272 4018 4346
rect 4214 4344 4470 4348
rect 5856 4346 5904 4422
rect 4214 4272 4472 4344
rect 4420 4270 4472 4272
rect 4928 4270 5186 4344
rect 5644 4272 5904 4346
rect 4930 4268 5186 4270
rect 1302 4162 2690 4224
rect 5968 4162 6168 4284
rect 1302 4024 1502 4162
rect 5734 4154 6168 4162
rect 5734 4118 5746 4154
rect 5788 4118 6168 4154
rect 5734 4112 6168 4118
rect 5968 4084 6168 4112
<< via1 >>
rect 2388 4588 2474 4682
rect 6178 4582 6272 4706
<< metal2 >>
rect 6178 4706 6272 4716
rect 2388 4688 2474 4692
rect 2388 4682 6178 4688
rect 2474 4606 6178 4682
rect 2388 4578 2474 4588
rect 6272 4606 6320 4688
rect 6178 4572 6272 4582
use sky130_fd_pr__pfet_01v8_BG9S83  sky130_fd_pr__pfet_01v8_BG9S83_0
timestamp 1708425308
transform 0 1 3353 -1 0 4916
box -226 -919 226 919
use sky130_fd_pr__pfet_01v8_6QP7WZ  XM1
timestamp 1707817411
transform 0 1 4985 -1 0 4916
box -226 -819 226 819
use sky130_fd_pr__nfet_01v8_8LLWK3  XM2
timestamp 1707817411
transform 0 1 4700 -1 0 4308
box -226 -410 226 410
use sky130_fd_pr__nfet_01v8_8LLWK3  XM3
timestamp 1707817411
transform 0 1 5414 -1 0 4308
box -226 -410 226 410
use sky130_fd_pr__pfet_01v8_SKJLLK  XM4
timestamp 0
transform 1 0 5997 0 1 5766
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_8YFQNF  XM5
timestamp 1707817411
transform 0 -1 4116 1 0 4308
box -226 -280 226 280
use sky130_fd_pr__pfet_01v8_GJYSVV  XM6
timestamp 1707817411
transform 0 1 2129 -1 0 4748
box -396 -319 396 319
use sky130_fd_pr__nfet_01v8_U4BYG2  XM7
timestamp 1707817411
transform 1 0 3148 0 1 4376
box -696 -310 696 310
use sky130_fd_pr__pfet_01v8_SKP3AN  XM8
timestamp 1707817411
transform 0 1 4065 1 0 5366
box -226 -2255 226 2255
<< labels >>
flabel metal1 1302 5410 1502 5610 0 FreeSans 256 0 0 0 vdd
port 3 nsew
flabel metal1 1302 4404 1502 4604 0 FreeSans 256 0 0 0 qa
port 0 nsew
flabel metal1 1302 4024 1502 4224 0 FreeSans 256 0 0 0 qb
port 1 nsew
flabel metal1 5968 4084 6168 4284 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 6124 4548 6324 4748 0 FreeSans 256 0 0 0 cp_out
port 2 nsew
flabel metal1 1298 4888 1498 5088 0 FreeSans 256 0 0 0 cp_bias
port 5 nsew
<< end >>
