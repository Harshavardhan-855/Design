magic
tech sky130A
magscale 1 2
timestamp 1706790953
<< error_p >>
rect -365 154 -307 160
rect -173 154 -115 160
rect 19 154 77 160
rect 211 154 269 160
rect 403 154 461 160
rect -365 120 -353 154
rect -173 120 -161 154
rect 19 120 31 154
rect 211 120 223 154
rect 403 120 415 154
rect -365 114 -307 120
rect -173 114 -115 120
rect 19 114 77 120
rect 211 114 269 120
rect 403 114 461 120
rect -461 -120 -403 -114
rect -269 -120 -211 -114
rect -77 -120 -19 -114
rect 115 -120 173 -114
rect 307 -120 365 -114
rect -461 -154 -449 -120
rect -269 -154 -257 -120
rect -77 -154 -65 -120
rect 115 -154 127 -120
rect 307 -154 319 -120
rect -461 -160 -403 -154
rect -269 -160 -211 -154
rect -77 -160 -19 -154
rect 115 -160 173 -154
rect 307 -160 365 -154
<< pwell >>
rect -647 -292 647 292
<< nmos >>
rect -447 -82 -417 82
rect -351 -82 -321 82
rect -255 -82 -225 82
rect -159 -82 -129 82
rect -63 -82 -33 82
rect 33 -82 63 82
rect 129 -82 159 82
rect 225 -82 255 82
rect 321 -82 351 82
rect 417 -82 447 82
<< ndiff >>
rect -509 70 -447 82
rect -509 -70 -497 70
rect -463 -70 -447 70
rect -509 -82 -447 -70
rect -417 70 -351 82
rect -417 -70 -401 70
rect -367 -70 -351 70
rect -417 -82 -351 -70
rect -321 70 -255 82
rect -321 -70 -305 70
rect -271 -70 -255 70
rect -321 -82 -255 -70
rect -225 70 -159 82
rect -225 -70 -209 70
rect -175 -70 -159 70
rect -225 -82 -159 -70
rect -129 70 -63 82
rect -129 -70 -113 70
rect -79 -70 -63 70
rect -129 -82 -63 -70
rect -33 70 33 82
rect -33 -70 -17 70
rect 17 -70 33 70
rect -33 -82 33 -70
rect 63 70 129 82
rect 63 -70 79 70
rect 113 -70 129 70
rect 63 -82 129 -70
rect 159 70 225 82
rect 159 -70 175 70
rect 209 -70 225 70
rect 159 -82 225 -70
rect 255 70 321 82
rect 255 -70 271 70
rect 305 -70 321 70
rect 255 -82 321 -70
rect 351 70 417 82
rect 351 -70 367 70
rect 401 -70 417 70
rect 351 -82 417 -70
rect 447 70 509 82
rect 447 -70 463 70
rect 497 -70 509 70
rect 447 -82 509 -70
<< ndiffc >>
rect -497 -70 -463 70
rect -401 -70 -367 70
rect -305 -70 -271 70
rect -209 -70 -175 70
rect -113 -70 -79 70
rect -17 -70 17 70
rect 79 -70 113 70
rect 175 -70 209 70
rect 271 -70 305 70
rect 367 -70 401 70
rect 463 -70 497 70
<< psubdiff >>
rect -611 222 -515 256
rect 515 222 611 256
rect -611 160 -577 222
rect 577 160 611 222
rect -611 -222 -577 -160
rect 577 -222 611 -160
rect -611 -256 -515 -222
rect 515 -256 611 -222
<< psubdiffcont >>
rect -515 222 515 256
rect -611 -160 -577 160
rect 577 -160 611 160
rect -515 -256 515 -222
<< poly >>
rect -369 154 -303 170
rect -369 120 -353 154
rect -319 120 -303 154
rect -447 82 -417 108
rect -369 104 -303 120
rect -177 154 -111 170
rect -177 120 -161 154
rect -127 120 -111 154
rect -351 82 -321 104
rect -255 82 -225 108
rect -177 104 -111 120
rect 15 154 81 170
rect 15 120 31 154
rect 65 120 81 154
rect -159 82 -129 104
rect -63 82 -33 108
rect 15 104 81 120
rect 207 154 273 170
rect 207 120 223 154
rect 257 120 273 154
rect 33 82 63 104
rect 129 82 159 108
rect 207 104 273 120
rect 399 154 465 170
rect 399 120 415 154
rect 449 120 465 154
rect 225 82 255 104
rect 321 82 351 108
rect 399 104 465 120
rect 417 82 447 104
rect -447 -104 -417 -82
rect -465 -120 -399 -104
rect -351 -108 -321 -82
rect -255 -104 -225 -82
rect -465 -154 -449 -120
rect -415 -154 -399 -120
rect -465 -170 -399 -154
rect -273 -120 -207 -104
rect -159 -108 -129 -82
rect -63 -104 -33 -82
rect -273 -154 -257 -120
rect -223 -154 -207 -120
rect -273 -170 -207 -154
rect -81 -120 -15 -104
rect 33 -108 63 -82
rect 129 -104 159 -82
rect -81 -154 -65 -120
rect -31 -154 -15 -120
rect -81 -170 -15 -154
rect 111 -120 177 -104
rect 225 -108 255 -82
rect 321 -104 351 -82
rect 111 -154 127 -120
rect 161 -154 177 -120
rect 111 -170 177 -154
rect 303 -120 369 -104
rect 417 -108 447 -82
rect 303 -154 319 -120
rect 353 -154 369 -120
rect 303 -170 369 -154
<< polycont >>
rect -353 120 -319 154
rect -161 120 -127 154
rect 31 120 65 154
rect 223 120 257 154
rect 415 120 449 154
rect -449 -154 -415 -120
rect -257 -154 -223 -120
rect -65 -154 -31 -120
rect 127 -154 161 -120
rect 319 -154 353 -120
<< locali >>
rect -611 222 -515 256
rect 515 222 611 256
rect -611 160 -577 222
rect 577 160 611 222
rect -369 120 -353 154
rect -319 120 -303 154
rect -177 120 -161 154
rect -127 120 -111 154
rect 15 120 31 154
rect 65 120 81 154
rect 207 120 223 154
rect 257 120 273 154
rect 399 120 415 154
rect 449 120 465 154
rect -497 70 -463 86
rect -497 -86 -463 -70
rect -401 70 -367 86
rect -401 -86 -367 -70
rect -305 70 -271 86
rect -305 -86 -271 -70
rect -209 70 -175 86
rect -209 -86 -175 -70
rect -113 70 -79 86
rect -113 -86 -79 -70
rect -17 70 17 86
rect -17 -86 17 -70
rect 79 70 113 86
rect 79 -86 113 -70
rect 175 70 209 86
rect 175 -86 209 -70
rect 271 70 305 86
rect 271 -86 305 -70
rect 367 70 401 86
rect 367 -86 401 -70
rect 463 70 497 86
rect 463 -86 497 -70
rect -465 -154 -449 -120
rect -415 -154 -399 -120
rect -273 -154 -257 -120
rect -223 -154 -207 -120
rect -81 -154 -65 -120
rect -31 -154 -15 -120
rect 111 -154 127 -120
rect 161 -154 177 -120
rect 303 -154 319 -120
rect 353 -154 369 -120
rect -611 -222 -577 -160
rect 577 -222 611 -160
rect -611 -256 -515 -222
rect 515 -256 611 -222
<< viali >>
rect -353 120 -319 154
rect -161 120 -127 154
rect 31 120 65 154
rect 223 120 257 154
rect 415 120 449 154
rect -497 -70 -463 70
rect -401 -70 -367 70
rect -305 -70 -271 70
rect -209 -70 -175 70
rect -113 -70 -79 70
rect -17 -70 17 70
rect 79 -70 113 70
rect 175 -70 209 70
rect 271 -70 305 70
rect 367 -70 401 70
rect 463 -70 497 70
rect -449 -154 -415 -120
rect -257 -154 -223 -120
rect -65 -154 -31 -120
rect 127 -154 161 -120
rect 319 -154 353 -120
<< metal1 >>
rect -365 154 -307 160
rect -365 120 -353 154
rect -319 120 -307 154
rect -365 114 -307 120
rect -173 154 -115 160
rect -173 120 -161 154
rect -127 120 -115 154
rect -173 114 -115 120
rect 19 154 77 160
rect 19 120 31 154
rect 65 120 77 154
rect 19 114 77 120
rect 211 154 269 160
rect 211 120 223 154
rect 257 120 269 154
rect 211 114 269 120
rect 403 154 461 160
rect 403 120 415 154
rect 449 120 461 154
rect 403 114 461 120
rect -503 70 -457 82
rect -503 -70 -497 70
rect -463 -70 -457 70
rect -503 -82 -457 -70
rect -407 70 -361 82
rect -407 -70 -401 70
rect -367 -70 -361 70
rect -407 -82 -361 -70
rect -311 70 -265 82
rect -311 -70 -305 70
rect -271 -70 -265 70
rect -311 -82 -265 -70
rect -215 70 -169 82
rect -215 -70 -209 70
rect -175 -70 -169 70
rect -215 -82 -169 -70
rect -119 70 -73 82
rect -119 -70 -113 70
rect -79 -70 -73 70
rect -119 -82 -73 -70
rect -23 70 23 82
rect -23 -70 -17 70
rect 17 -70 23 70
rect -23 -82 23 -70
rect 73 70 119 82
rect 73 -70 79 70
rect 113 -70 119 70
rect 73 -82 119 -70
rect 169 70 215 82
rect 169 -70 175 70
rect 209 -70 215 70
rect 169 -82 215 -70
rect 265 70 311 82
rect 265 -70 271 70
rect 305 -70 311 70
rect 265 -82 311 -70
rect 361 70 407 82
rect 361 -70 367 70
rect 401 -70 407 70
rect 361 -82 407 -70
rect 457 70 503 82
rect 457 -70 463 70
rect 497 -70 503 70
rect 457 -82 503 -70
rect -461 -120 -403 -114
rect -461 -154 -449 -120
rect -415 -154 -403 -120
rect -461 -160 -403 -154
rect -269 -120 -211 -114
rect -269 -154 -257 -120
rect -223 -154 -211 -120
rect -269 -160 -211 -154
rect -77 -120 -19 -114
rect -77 -154 -65 -120
rect -31 -154 -19 -120
rect -77 -160 -19 -154
rect 115 -120 173 -114
rect 115 -154 127 -120
rect 161 -154 173 -120
rect 115 -160 173 -154
rect 307 -120 365 -114
rect 307 -154 319 -120
rect 353 -154 365 -120
rect 307 -160 365 -154
<< properties >>
string FIXED_BBOX -594 -239 594 239
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.820 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
