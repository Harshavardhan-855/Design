magic
tech sky130A
magscale 1 2
timestamp 1709561889
<< error_p >>
rect -29 142 29 148
rect -29 108 -17 142
rect -29 102 29 108
rect -29 -108 29 -102
rect -29 -142 -17 -108
rect -29 -148 29 -142
<< pwell >>
rect -226 -280 226 280
<< nmos >>
rect -30 -70 30 70
<< ndiff >>
rect -88 58 -30 70
rect -88 -58 -76 58
rect -42 -58 -30 58
rect -88 -70 -30 -58
rect 30 58 88 70
rect 30 -58 42 58
rect 76 -58 88 58
rect 30 -70 88 -58
<< ndiffc >>
rect -76 -58 -42 58
rect 42 -58 76 58
<< psubdiff >>
rect -190 210 -94 244
rect 94 210 190 244
rect -190 148 -156 210
rect 156 148 190 210
rect -190 -210 -156 -148
rect 156 -210 190 -148
rect -190 -244 -94 -210
rect 94 -244 190 -210
<< psubdiffcont >>
rect -94 210 94 244
rect -190 -148 -156 148
rect 156 -148 190 148
rect -94 -244 94 -210
<< poly >>
rect -33 142 33 158
rect -33 108 -17 142
rect 17 108 33 142
rect -33 92 33 108
rect -30 70 30 92
rect -30 -92 30 -70
rect -33 -108 33 -92
rect -33 -142 -17 -108
rect 17 -142 33 -108
rect -33 -158 33 -142
<< polycont >>
rect -17 108 17 142
rect -17 -142 17 -108
<< locali >>
rect -190 210 -94 244
rect 94 210 190 244
rect -190 148 -156 210
rect 156 148 190 210
rect -33 108 -17 142
rect 17 108 33 142
rect -76 58 -42 74
rect -76 -74 -42 -58
rect 42 58 76 74
rect 42 -74 76 -58
rect -33 -142 -17 -108
rect 17 -142 33 -108
rect -190 -210 -156 -148
rect 156 -210 190 -148
rect -190 -244 -94 -210
rect 94 -244 190 -210
<< viali >>
rect -17 108 17 142
rect -76 -58 -42 58
rect 42 -58 76 58
rect -17 -142 17 -108
<< metal1 >>
rect -29 142 29 148
rect -29 108 -17 142
rect 17 108 29 142
rect -29 102 29 108
rect -82 58 -36 70
rect -82 -58 -76 58
rect -42 -58 -36 58
rect -82 -70 -36 -58
rect 36 58 82 70
rect 36 -58 42 58
rect 76 -58 82 58
rect 36 -70 82 -58
rect -29 -108 29 -102
rect -29 -142 -17 -108
rect 17 -142 29 -108
rect -29 -148 29 -142
<< properties >>
string FIXED_BBOX -173 -227 173 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
