magic
tech sky130A
magscale 1 2
timestamp 1706794580
<< pwell >>
rect -266 -846 266 846
<< psubdiff >>
rect -230 776 -134 810
rect 134 776 230 810
rect -230 714 -196 776
rect 196 714 230 776
rect -230 -776 -196 -714
rect 196 -776 230 -714
rect -230 -810 -134 -776
rect 134 -810 230 -776
<< psubdiffcont >>
rect -134 776 134 810
rect -230 -714 -196 714
rect 196 -714 230 714
rect -134 -810 134 -776
<< poly >>
rect -100 664 100 680
rect -100 630 -84 664
rect 84 630 100 664
rect -100 250 100 630
rect -100 -630 100 -250
rect -100 -664 -84 -630
rect 84 -664 100 -630
rect -100 -680 100 -664
<< polycont >>
rect -84 630 84 664
rect -84 -664 84 -630
<< npolyres >>
rect -100 -250 100 250
<< locali >>
rect -230 776 -134 810
rect 134 776 230 810
rect -230 714 -196 776
rect 196 714 230 776
rect -100 630 -84 664
rect 84 630 100 664
rect -100 -664 -84 -630
rect 84 -664 100 -630
rect -230 -776 -196 -714
rect 196 -776 230 -714
rect -230 -810 -134 -776
rect 134 -810 230 -776
<< viali >>
rect -84 630 84 664
rect -84 267 84 630
rect -84 -630 84 -267
rect -84 -664 84 -630
<< metal1 >>
rect -90 664 90 676
rect -90 267 -84 664
rect 84 267 90 664
rect -90 255 90 267
rect -90 -267 90 -255
rect -90 -664 -84 -267
rect 84 -664 90 -267
rect -90 -676 90 -664
<< properties >>
string FIXED_BBOX -213 -793 213 793
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 1.0 l 2.5 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 120.5 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
