magic
tech sky130A
magscale 1 2
timestamp 1709130382
<< error_p >>
rect -1037 123 -979 129
rect -845 123 -787 129
rect -653 123 -595 129
rect -461 123 -403 129
rect -269 123 -211 129
rect -77 123 -19 129
rect 115 123 173 129
rect 307 123 365 129
rect 499 123 557 129
rect 691 123 749 129
rect 883 123 941 129
rect 1075 123 1133 129
rect -1037 89 -1025 123
rect -845 89 -833 123
rect -653 89 -641 123
rect -461 89 -449 123
rect -269 89 -257 123
rect -77 89 -65 123
rect 115 89 127 123
rect 307 89 319 123
rect 499 89 511 123
rect 691 89 703 123
rect 883 89 895 123
rect 1075 89 1087 123
rect -1037 83 -979 89
rect -845 83 -787 89
rect -653 83 -595 89
rect -461 83 -403 89
rect -269 83 -211 89
rect -77 83 -19 89
rect 115 83 173 89
rect 307 83 365 89
rect 499 83 557 89
rect 691 83 749 89
rect 883 83 941 89
rect 1075 83 1133 89
rect -1133 -89 -1075 -83
rect -941 -89 -883 -83
rect -749 -89 -691 -83
rect -557 -89 -499 -83
rect -365 -89 -307 -83
rect -173 -89 -115 -83
rect 19 -89 77 -83
rect 211 -89 269 -83
rect 403 -89 461 -83
rect 595 -89 653 -83
rect 787 -89 845 -83
rect 979 -89 1037 -83
rect -1133 -123 -1121 -89
rect -941 -123 -929 -89
rect -749 -123 -737 -89
rect -557 -123 -545 -89
rect -365 -123 -353 -89
rect -173 -123 -161 -89
rect 19 -123 31 -89
rect 211 -123 223 -89
rect 403 -123 415 -89
rect 595 -123 607 -89
rect 787 -123 799 -89
rect 979 -123 991 -89
rect -1133 -129 -1075 -123
rect -941 -129 -883 -123
rect -749 -129 -691 -123
rect -557 -129 -499 -123
rect -365 -129 -307 -123
rect -173 -129 -115 -123
rect 19 -129 77 -123
rect 211 -129 269 -123
rect 403 -129 461 -123
rect 595 -129 653 -123
rect 787 -129 845 -123
rect 979 -129 1037 -123
<< nwell >>
rect -1319 -261 1319 261
<< pmos >>
rect -1119 -42 -1089 42
rect -1023 -42 -993 42
rect -927 -42 -897 42
rect -831 -42 -801 42
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
rect 801 -42 831 42
rect 897 -42 927 42
rect 993 -42 1023 42
rect 1089 -42 1119 42
<< pdiff >>
rect -1181 30 -1119 42
rect -1181 -30 -1169 30
rect -1135 -30 -1119 30
rect -1181 -42 -1119 -30
rect -1089 30 -1023 42
rect -1089 -30 -1073 30
rect -1039 -30 -1023 30
rect -1089 -42 -1023 -30
rect -993 30 -927 42
rect -993 -30 -977 30
rect -943 -30 -927 30
rect -993 -42 -927 -30
rect -897 30 -831 42
rect -897 -30 -881 30
rect -847 -30 -831 30
rect -897 -42 -831 -30
rect -801 30 -735 42
rect -801 -30 -785 30
rect -751 -30 -735 30
rect -801 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 801 42
rect 735 -30 751 30
rect 785 -30 801 30
rect 735 -42 801 -30
rect 831 30 897 42
rect 831 -30 847 30
rect 881 -30 897 30
rect 831 -42 897 -30
rect 927 30 993 42
rect 927 -30 943 30
rect 977 -30 993 30
rect 927 -42 993 -30
rect 1023 30 1089 42
rect 1023 -30 1039 30
rect 1073 -30 1089 30
rect 1023 -42 1089 -30
rect 1119 30 1181 42
rect 1119 -30 1135 30
rect 1169 -30 1181 30
rect 1119 -42 1181 -30
<< pdiffc >>
rect -1169 -30 -1135 30
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect 1135 -30 1169 30
<< nsubdiff >>
rect -1283 191 -1187 225
rect 1187 191 1283 225
rect -1283 129 -1249 191
rect 1249 129 1283 191
rect -1283 -191 -1249 -129
rect 1249 -191 1283 -129
rect -1283 -225 -1187 -191
rect 1187 -225 1283 -191
<< nsubdiffcont >>
rect -1187 191 1187 225
rect -1283 -129 -1249 129
rect 1249 -129 1283 129
rect -1187 -225 1187 -191
<< poly >>
rect -1041 123 -975 139
rect -1041 89 -1025 123
rect -991 89 -975 123
rect -1041 73 -975 89
rect -849 123 -783 139
rect -849 89 -833 123
rect -799 89 -783 123
rect -849 73 -783 89
rect -657 123 -591 139
rect -657 89 -641 123
rect -607 89 -591 123
rect -657 73 -591 89
rect -465 123 -399 139
rect -465 89 -449 123
rect -415 89 -399 123
rect -465 73 -399 89
rect -273 123 -207 139
rect -273 89 -257 123
rect -223 89 -207 123
rect -273 73 -207 89
rect -81 123 -15 139
rect -81 89 -65 123
rect -31 89 -15 123
rect -81 73 -15 89
rect 111 123 177 139
rect 111 89 127 123
rect 161 89 177 123
rect 111 73 177 89
rect 303 123 369 139
rect 303 89 319 123
rect 353 89 369 123
rect 303 73 369 89
rect 495 123 561 139
rect 495 89 511 123
rect 545 89 561 123
rect 495 73 561 89
rect 687 123 753 139
rect 687 89 703 123
rect 737 89 753 123
rect 687 73 753 89
rect 879 123 945 139
rect 879 89 895 123
rect 929 89 945 123
rect 879 73 945 89
rect 1071 123 1137 139
rect 1071 89 1087 123
rect 1121 89 1137 123
rect 1071 73 1137 89
rect -1119 42 -1089 68
rect -1023 42 -993 73
rect -927 42 -897 68
rect -831 42 -801 73
rect -735 42 -705 68
rect -639 42 -609 73
rect -543 42 -513 68
rect -447 42 -417 73
rect -351 42 -321 68
rect -255 42 -225 73
rect -159 42 -129 68
rect -63 42 -33 73
rect 33 42 63 68
rect 129 42 159 73
rect 225 42 255 68
rect 321 42 351 73
rect 417 42 447 68
rect 513 42 543 73
rect 609 42 639 68
rect 705 42 735 73
rect 801 42 831 68
rect 897 42 927 73
rect 993 42 1023 68
rect 1089 42 1119 73
rect -1119 -73 -1089 -42
rect -1023 -68 -993 -42
rect -927 -73 -897 -42
rect -831 -68 -801 -42
rect -735 -73 -705 -42
rect -639 -68 -609 -42
rect -543 -73 -513 -42
rect -447 -68 -417 -42
rect -351 -73 -321 -42
rect -255 -68 -225 -42
rect -159 -73 -129 -42
rect -63 -68 -33 -42
rect 33 -73 63 -42
rect 129 -68 159 -42
rect 225 -73 255 -42
rect 321 -68 351 -42
rect 417 -73 447 -42
rect 513 -68 543 -42
rect 609 -73 639 -42
rect 705 -68 735 -42
rect 801 -73 831 -42
rect 897 -68 927 -42
rect 993 -73 1023 -42
rect 1089 -68 1119 -42
rect -1137 -89 -1071 -73
rect -1137 -123 -1121 -89
rect -1087 -123 -1071 -89
rect -1137 -139 -1071 -123
rect -945 -89 -879 -73
rect -945 -123 -929 -89
rect -895 -123 -879 -89
rect -945 -139 -879 -123
rect -753 -89 -687 -73
rect -753 -123 -737 -89
rect -703 -123 -687 -89
rect -753 -139 -687 -123
rect -561 -89 -495 -73
rect -561 -123 -545 -89
rect -511 -123 -495 -89
rect -561 -139 -495 -123
rect -369 -89 -303 -73
rect -369 -123 -353 -89
rect -319 -123 -303 -89
rect -369 -139 -303 -123
rect -177 -89 -111 -73
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect -177 -139 -111 -123
rect 15 -89 81 -73
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 15 -139 81 -123
rect 207 -89 273 -73
rect 207 -123 223 -89
rect 257 -123 273 -89
rect 207 -139 273 -123
rect 399 -89 465 -73
rect 399 -123 415 -89
rect 449 -123 465 -89
rect 399 -139 465 -123
rect 591 -89 657 -73
rect 591 -123 607 -89
rect 641 -123 657 -89
rect 591 -139 657 -123
rect 783 -89 849 -73
rect 783 -123 799 -89
rect 833 -123 849 -89
rect 783 -139 849 -123
rect 975 -89 1041 -73
rect 975 -123 991 -89
rect 1025 -123 1041 -89
rect 975 -139 1041 -123
<< polycont >>
rect -1025 89 -991 123
rect -833 89 -799 123
rect -641 89 -607 123
rect -449 89 -415 123
rect -257 89 -223 123
rect -65 89 -31 123
rect 127 89 161 123
rect 319 89 353 123
rect 511 89 545 123
rect 703 89 737 123
rect 895 89 929 123
rect 1087 89 1121 123
rect -1121 -123 -1087 -89
rect -929 -123 -895 -89
rect -737 -123 -703 -89
rect -545 -123 -511 -89
rect -353 -123 -319 -89
rect -161 -123 -127 -89
rect 31 -123 65 -89
rect 223 -123 257 -89
rect 415 -123 449 -89
rect 607 -123 641 -89
rect 799 -123 833 -89
rect 991 -123 1025 -89
<< locali >>
rect -1283 191 -1187 225
rect 1187 191 1283 225
rect -1283 129 -1249 191
rect 1249 129 1283 191
rect -1041 89 -1025 123
rect -991 89 -975 123
rect -849 89 -833 123
rect -799 89 -783 123
rect -657 89 -641 123
rect -607 89 -591 123
rect -465 89 -449 123
rect -415 89 -399 123
rect -273 89 -257 123
rect -223 89 -207 123
rect -81 89 -65 123
rect -31 89 -15 123
rect 111 89 127 123
rect 161 89 177 123
rect 303 89 319 123
rect 353 89 369 123
rect 495 89 511 123
rect 545 89 561 123
rect 687 89 703 123
rect 737 89 753 123
rect 879 89 895 123
rect 929 89 945 123
rect 1071 89 1087 123
rect 1121 89 1137 123
rect -1169 30 -1135 46
rect -1169 -46 -1135 -30
rect -1073 30 -1039 46
rect -1073 -46 -1039 -30
rect -977 30 -943 46
rect -977 -46 -943 -30
rect -881 30 -847 46
rect -881 -46 -847 -30
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect 847 30 881 46
rect 847 -46 881 -30
rect 943 30 977 46
rect 943 -46 977 -30
rect 1039 30 1073 46
rect 1039 -46 1073 -30
rect 1135 30 1169 46
rect 1135 -46 1169 -30
rect -1137 -123 -1121 -89
rect -1087 -123 -1071 -89
rect -945 -123 -929 -89
rect -895 -123 -879 -89
rect -753 -123 -737 -89
rect -703 -123 -687 -89
rect -561 -123 -545 -89
rect -511 -123 -495 -89
rect -369 -123 -353 -89
rect -319 -123 -303 -89
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 207 -123 223 -89
rect 257 -123 273 -89
rect 399 -123 415 -89
rect 449 -123 465 -89
rect 591 -123 607 -89
rect 641 -123 657 -89
rect 783 -123 799 -89
rect 833 -123 849 -89
rect 975 -123 991 -89
rect 1025 -123 1041 -89
rect -1283 -191 -1249 -129
rect 1249 -191 1283 -129
rect -1283 -225 -1187 -191
rect 1187 -225 1283 -191
<< viali >>
rect -1025 89 -991 123
rect -833 89 -799 123
rect -641 89 -607 123
rect -449 89 -415 123
rect -257 89 -223 123
rect -65 89 -31 123
rect 127 89 161 123
rect 319 89 353 123
rect 511 89 545 123
rect 703 89 737 123
rect 895 89 929 123
rect 1087 89 1121 123
rect -1169 -30 -1135 30
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect 1135 -30 1169 30
rect -1121 -123 -1087 -89
rect -929 -123 -895 -89
rect -737 -123 -703 -89
rect -545 -123 -511 -89
rect -353 -123 -319 -89
rect -161 -123 -127 -89
rect 31 -123 65 -89
rect 223 -123 257 -89
rect 415 -123 449 -89
rect 607 -123 641 -89
rect 799 -123 833 -89
rect 991 -123 1025 -89
<< metal1 >>
rect -1037 123 -979 129
rect -1037 89 -1025 123
rect -991 89 -979 123
rect -1037 83 -979 89
rect -845 123 -787 129
rect -845 89 -833 123
rect -799 89 -787 123
rect -845 83 -787 89
rect -653 123 -595 129
rect -653 89 -641 123
rect -607 89 -595 123
rect -653 83 -595 89
rect -461 123 -403 129
rect -461 89 -449 123
rect -415 89 -403 123
rect -461 83 -403 89
rect -269 123 -211 129
rect -269 89 -257 123
rect -223 89 -211 123
rect -269 83 -211 89
rect -77 123 -19 129
rect -77 89 -65 123
rect -31 89 -19 123
rect -77 83 -19 89
rect 115 123 173 129
rect 115 89 127 123
rect 161 89 173 123
rect 115 83 173 89
rect 307 123 365 129
rect 307 89 319 123
rect 353 89 365 123
rect 307 83 365 89
rect 499 123 557 129
rect 499 89 511 123
rect 545 89 557 123
rect 499 83 557 89
rect 691 123 749 129
rect 691 89 703 123
rect 737 89 749 123
rect 691 83 749 89
rect 883 123 941 129
rect 883 89 895 123
rect 929 89 941 123
rect 883 83 941 89
rect 1075 123 1133 129
rect 1075 89 1087 123
rect 1121 89 1133 123
rect 1075 83 1133 89
rect -1175 30 -1129 42
rect -1175 -30 -1169 30
rect -1135 -30 -1129 30
rect -1175 -42 -1129 -30
rect -1079 30 -1033 42
rect -1079 -30 -1073 30
rect -1039 -30 -1033 30
rect -1079 -42 -1033 -30
rect -983 30 -937 42
rect -983 -30 -977 30
rect -943 -30 -937 30
rect -983 -42 -937 -30
rect -887 30 -841 42
rect -887 -30 -881 30
rect -847 -30 -841 30
rect -887 -42 -841 -30
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
rect 841 30 887 42
rect 841 -30 847 30
rect 881 -30 887 30
rect 841 -42 887 -30
rect 937 30 983 42
rect 937 -30 943 30
rect 977 -30 983 30
rect 937 -42 983 -30
rect 1033 30 1079 42
rect 1033 -30 1039 30
rect 1073 -30 1079 30
rect 1033 -42 1079 -30
rect 1129 30 1175 42
rect 1129 -30 1135 30
rect 1169 -30 1175 30
rect 1129 -42 1175 -30
rect -1133 -89 -1075 -83
rect -1133 -123 -1121 -89
rect -1087 -123 -1075 -89
rect -1133 -129 -1075 -123
rect -941 -89 -883 -83
rect -941 -123 -929 -89
rect -895 -123 -883 -89
rect -941 -129 -883 -123
rect -749 -89 -691 -83
rect -749 -123 -737 -89
rect -703 -123 -691 -89
rect -749 -129 -691 -123
rect -557 -89 -499 -83
rect -557 -123 -545 -89
rect -511 -123 -499 -89
rect -557 -129 -499 -123
rect -365 -89 -307 -83
rect -365 -123 -353 -89
rect -319 -123 -307 -89
rect -365 -129 -307 -123
rect -173 -89 -115 -83
rect -173 -123 -161 -89
rect -127 -123 -115 -89
rect -173 -129 -115 -123
rect 19 -89 77 -83
rect 19 -123 31 -89
rect 65 -123 77 -89
rect 19 -129 77 -123
rect 211 -89 269 -83
rect 211 -123 223 -89
rect 257 -123 269 -89
rect 211 -129 269 -123
rect 403 -89 461 -83
rect 403 -123 415 -89
rect 449 -123 461 -89
rect 403 -129 461 -123
rect 595 -89 653 -83
rect 595 -123 607 -89
rect 641 -123 653 -89
rect 595 -129 653 -123
rect 787 -89 845 -83
rect 787 -123 799 -89
rect 833 -123 845 -89
rect 787 -129 845 -123
rect 979 -89 1037 -83
rect 979 -123 991 -89
rect 1025 -123 1037 -89
rect 979 -129 1037 -123
<< properties >>
string FIXED_BBOX -1266 -208 1266 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
