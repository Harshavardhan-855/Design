** sch_path: /home/harsh/design/xschem/untitledppp.sch
**.subckt untitledppp
x1 net1 net2 net3 net4 net5 net6 pfd
x2 net7 net8 net9 net10 net11 net12 cp_schem
**.ends

* expanding   symbol:  PLL_FOLDER/pfd.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/pfd.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/pfd.sch
.subckt pfd VSS VDD A QA QB B
*.iopin VDD
*.iopin A
*.iopin B
*.iopin QA
*.iopin QB
*.iopin VSS
x1 A VDD reset VSS VSS VDD VDD QA net2 sky130_fd_sc_hd__dfrbp_2
x2 QA QB VSS VSS VDD VDD net1 sky130_fd_sc_hd__and2_2
x3 B VDD reset VSS VSS VDD VDD QB net3 sky130_fd_sc_hd__dfrbp_2
x4 net1 VSS VSS VDD VDD reset sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  PLL_FOLDER/cp/cp_schem.sym # of pins=6
** sym_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sym
** sch_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sch
.subckt cp_schem vdd cp_bias qa cp_out qb vss
*.ipin qa
*.ipin qb
*.opin cp_out
*.iopin vdd
*.iopin vss
*.ipin cp_bias
XM1 n1 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 n1 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 bias bias vss vss sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 n2 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 n3 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 cp_out qa n2 vdd sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 cp_out qb n3 vss sky130_fd_pr__nfet_01v8 L=5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 bias cp_bias vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
.ends

.end
